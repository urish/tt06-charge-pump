magic
tech sky130A
magscale 1 2
timestamp 1711870259
<< nwell >>
rect -241 -369 241 369
<< pmos >>
rect -45 -150 45 150
<< pdiff >>
rect -103 138 -45 150
rect -103 -138 -91 138
rect -57 -138 -45 138
rect -103 -150 -45 -138
rect 45 138 103 150
rect 45 -138 57 138
rect 91 -138 103 138
rect 45 -150 103 -138
<< pdiffc >>
rect -91 -138 -57 138
rect 57 -138 91 138
<< nsubdiff >>
rect -205 299 -109 333
rect 109 299 205 333
rect -205 237 -171 299
rect 171 237 205 299
rect -205 -299 -171 -237
rect 171 -299 205 -237
rect -205 -333 -109 -299
rect 109 -333 205 -299
<< nsubdiffcont >>
rect -109 299 109 333
rect -205 -237 -171 237
rect 171 -237 205 237
rect -109 -333 109 -299
<< poly >>
rect -45 231 45 247
rect -45 197 -29 231
rect 29 197 45 231
rect -45 150 45 197
rect -45 -197 45 -150
rect -45 -231 -29 -197
rect 29 -231 45 -197
rect -45 -247 45 -231
<< polycont >>
rect -29 197 29 231
rect -29 -231 29 -197
<< locali >>
rect -205 299 -109 333
rect 109 299 205 333
rect -205 237 -171 299
rect 171 237 205 299
rect -45 197 -29 231
rect 29 197 45 231
rect -91 138 -57 154
rect -91 -154 -57 -138
rect 57 138 91 154
rect 57 -154 91 -138
rect -45 -231 -29 -197
rect 29 -231 45 -197
rect -205 -299 -171 -237
rect 171 -299 205 -237
rect -205 -333 -109 -299
rect 109 -333 205 -299
<< viali >>
rect -29 197 29 231
rect -91 -138 -57 138
rect 57 -138 91 138
rect -29 -231 29 -197
<< metal1 >>
rect -41 231 41 237
rect -41 197 -29 231
rect 29 197 41 231
rect -41 191 41 197
rect -97 138 -51 150
rect -97 -138 -91 138
rect -57 -138 -51 138
rect -97 -150 -51 -138
rect 51 138 97 150
rect 51 -138 57 138
rect 91 -138 97 138
rect 51 -150 97 -138
rect -41 -197 41 -191
rect -41 -231 -29 -197
rect 29 -231 41 -197
rect -41 -237 41 -231
<< properties >>
string FIXED_BBOX -188 -316 188 316
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.45 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
