magic
tech sky130A
timestamp 1711870259
<< pwell >>
rect -2134 -2668 2134 2668
<< psubdiff >>
rect -2116 2633 -2068 2650
rect 2068 2633 2116 2650
rect -2116 2602 -2099 2633
rect 2099 2602 2116 2633
rect -2116 -2633 -2099 -2602
rect 2099 -2633 2116 -2602
rect -2116 -2650 -2068 -2633
rect 2068 -2650 2116 -2633
<< psubdiffcont >>
rect -2068 2633 2068 2650
rect -2116 -2602 -2099 2602
rect 2099 -2602 2116 2602
rect -2068 -2650 2068 -2633
<< xpolycontact >>
rect -2051 -2585 -2016 -2369
rect 2016 -2585 2051 -2369
<< xpolyres >>
rect -2051 2550 -1933 2585
rect -2051 -2369 -2016 2550
rect -1968 -2282 -1933 2550
rect -1885 2550 -1767 2585
rect -1885 -2282 -1850 2550
rect -1968 -2317 -1850 -2282
rect -1802 -2282 -1767 2550
rect -1719 2550 -1601 2585
rect -1719 -2282 -1684 2550
rect -1802 -2317 -1684 -2282
rect -1636 -2282 -1601 2550
rect -1553 2550 -1435 2585
rect -1553 -2282 -1518 2550
rect -1636 -2317 -1518 -2282
rect -1470 -2282 -1435 2550
rect -1387 2550 -1269 2585
rect -1387 -2282 -1352 2550
rect -1470 -2317 -1352 -2282
rect -1304 -2282 -1269 2550
rect -1221 2550 -1103 2585
rect -1221 -2282 -1186 2550
rect -1304 -2317 -1186 -2282
rect -1138 -2282 -1103 2550
rect -1055 2550 -937 2585
rect -1055 -2282 -1020 2550
rect -1138 -2317 -1020 -2282
rect -972 -2282 -937 2550
rect -889 2550 -771 2585
rect -889 -2282 -854 2550
rect -972 -2317 -854 -2282
rect -806 -2282 -771 2550
rect -723 2550 -605 2585
rect -723 -2282 -688 2550
rect -806 -2317 -688 -2282
rect -640 -2282 -605 2550
rect -557 2550 -439 2585
rect -557 -2282 -522 2550
rect -640 -2317 -522 -2282
rect -474 -2282 -439 2550
rect -391 2550 -273 2585
rect -391 -2282 -356 2550
rect -474 -2317 -356 -2282
rect -308 -2282 -273 2550
rect -225 2550 -107 2585
rect -225 -2282 -190 2550
rect -308 -2317 -190 -2282
rect -142 -2282 -107 2550
rect -59 2550 59 2585
rect -59 -2282 -24 2550
rect -142 -2317 -24 -2282
rect 24 -2282 59 2550
rect 107 2550 225 2585
rect 107 -2282 142 2550
rect 24 -2317 142 -2282
rect 190 -2282 225 2550
rect 273 2550 391 2585
rect 273 -2282 308 2550
rect 190 -2317 308 -2282
rect 356 -2282 391 2550
rect 439 2550 557 2585
rect 439 -2282 474 2550
rect 356 -2317 474 -2282
rect 522 -2282 557 2550
rect 605 2550 723 2585
rect 605 -2282 640 2550
rect 522 -2317 640 -2282
rect 688 -2282 723 2550
rect 771 2550 889 2585
rect 771 -2282 806 2550
rect 688 -2317 806 -2282
rect 854 -2282 889 2550
rect 937 2550 1055 2585
rect 937 -2282 972 2550
rect 854 -2317 972 -2282
rect 1020 -2282 1055 2550
rect 1103 2550 1221 2585
rect 1103 -2282 1138 2550
rect 1020 -2317 1138 -2282
rect 1186 -2282 1221 2550
rect 1269 2550 1387 2585
rect 1269 -2282 1304 2550
rect 1186 -2317 1304 -2282
rect 1352 -2282 1387 2550
rect 1435 2550 1553 2585
rect 1435 -2282 1470 2550
rect 1352 -2317 1470 -2282
rect 1518 -2282 1553 2550
rect 1601 2550 1719 2585
rect 1601 -2282 1636 2550
rect 1518 -2317 1636 -2282
rect 1684 -2282 1719 2550
rect 1767 2550 1885 2585
rect 1767 -2282 1802 2550
rect 1684 -2317 1802 -2282
rect 1850 -2282 1885 2550
rect 1933 2550 2051 2585
rect 1933 -2282 1968 2550
rect 1850 -2317 1968 -2282
rect 2016 -2369 2051 2550
<< locali >>
rect -2116 2633 -2068 2650
rect 2068 2633 2116 2650
rect -2116 2602 -2099 2633
rect 2099 2602 2116 2633
rect -2116 -2633 -2099 -2602
rect 2099 -2633 2116 -2602
rect -2116 -2650 -2068 -2633
rect 2068 -2650 2116 -2633
<< properties >>
string FIXED_BBOX -2107 -2641 2107 2641
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 49.02 m 1 nx 50 wmin 0.350 lmin 0.50 rho 2000 val 14.104meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
