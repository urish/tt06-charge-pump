VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_charge_pump
  CLASS BLOCK ;
  FOREIGN tt_um_urish_charge_pump ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 151.000 219.500 153.410 223.190 ;
        RECT 155.000 219.500 157.410 223.190 ;
      LAYER pwell ;
        RECT 151.000 216.000 153.410 219.100 ;
        RECT 155.000 216.000 157.410 219.100 ;
        RECT 148.000 189.500 157.960 198.600 ;
        RECT 149.500 160.500 159.460 169.600 ;
        RECT 150.500 119.500 160.460 128.600 ;
        RECT 150.000 78.000 159.960 87.100 ;
        RECT 106.550 7.550 149.230 60.910 ;
        RECT 149.650 7.550 154.980 63.770 ;
      LAYER li1 ;
        RECT 151.180 222.840 153.230 223.010 ;
        RECT 151.180 219.850 151.350 222.840 ;
        RECT 151.980 222.330 152.430 222.500 ;
        RECT 151.750 220.575 151.920 222.115 ;
        RECT 152.490 220.575 152.660 222.115 ;
        RECT 151.980 220.190 152.430 220.360 ;
        RECT 153.060 219.850 153.230 222.840 ;
        RECT 151.180 219.680 153.230 219.850 ;
        RECT 155.180 222.840 157.230 223.010 ;
        RECT 155.180 219.850 155.350 222.840 ;
        RECT 155.980 222.330 156.430 222.500 ;
        RECT 155.750 220.575 155.920 222.115 ;
        RECT 156.490 220.575 156.660 222.115 ;
        RECT 155.980 220.190 156.430 220.360 ;
        RECT 157.060 219.850 157.230 222.840 ;
        RECT 155.180 219.680 157.230 219.850 ;
        RECT 151.180 218.750 153.230 218.920 ;
        RECT 151.180 216.350 151.350 218.750 ;
        RECT 151.980 218.240 152.430 218.410 ;
        RECT 151.750 217.030 151.920 218.070 ;
        RECT 152.490 217.030 152.660 218.070 ;
        RECT 151.980 216.690 152.430 216.860 ;
        RECT 153.060 216.350 153.230 218.750 ;
        RECT 151.180 216.180 153.230 216.350 ;
        RECT 155.180 218.750 157.230 218.920 ;
        RECT 155.180 216.350 155.350 218.750 ;
        RECT 155.980 218.240 156.430 218.410 ;
        RECT 155.750 217.030 155.920 218.070 ;
        RECT 156.490 217.030 156.660 218.070 ;
        RECT 155.980 216.690 156.430 216.860 ;
        RECT 157.060 216.350 157.230 218.750 ;
        RECT 155.180 216.180 157.230 216.350 ;
        RECT 148.180 198.250 157.780 198.420 ;
        RECT 148.180 189.850 148.350 198.250 ;
        RECT 148.980 197.740 156.980 197.910 ;
        RECT 148.750 190.530 148.920 197.570 ;
        RECT 157.040 190.530 157.210 197.570 ;
        RECT 148.980 190.190 156.980 190.360 ;
        RECT 157.610 189.850 157.780 198.250 ;
        RECT 148.180 189.680 157.780 189.850 ;
        RECT 149.680 169.250 159.280 169.420 ;
        RECT 149.680 160.850 149.850 169.250 ;
        RECT 150.480 168.740 158.480 168.910 ;
        RECT 150.250 161.530 150.420 168.570 ;
        RECT 158.540 161.530 158.710 168.570 ;
        RECT 150.480 161.190 158.480 161.360 ;
        RECT 159.110 160.850 159.280 169.250 ;
        RECT 149.680 160.680 159.280 160.850 ;
        RECT 150.680 128.250 160.280 128.420 ;
        RECT 150.680 119.850 150.850 128.250 ;
        RECT 151.480 127.740 159.480 127.910 ;
        RECT 151.250 120.530 151.420 127.570 ;
        RECT 159.540 120.530 159.710 127.570 ;
        RECT 151.480 120.190 159.480 120.360 ;
        RECT 160.110 119.850 160.280 128.250 ;
        RECT 150.680 119.680 160.280 119.850 ;
        RECT 150.180 86.750 159.780 86.920 ;
        RECT 150.180 78.350 150.350 86.750 ;
        RECT 150.980 86.240 158.980 86.410 ;
        RECT 150.750 79.030 150.920 86.070 ;
        RECT 159.040 79.030 159.210 86.070 ;
        RECT 150.980 78.690 158.980 78.860 ;
        RECT 159.610 78.350 159.780 86.750 ;
        RECT 150.180 78.180 159.780 78.350 ;
        RECT 149.830 63.420 154.800 63.590 ;
        RECT 106.730 60.560 149.050 60.730 ;
        RECT 106.730 7.900 106.900 60.560 ;
        RECT 107.380 8.380 107.730 10.540 ;
        RECT 148.050 8.380 148.400 10.540 ;
        RECT 148.880 7.900 149.050 60.560 ;
        RECT 106.730 7.730 149.050 7.900 ;
        RECT 149.830 7.900 150.000 63.420 ;
        RECT 153.800 60.780 154.150 62.940 ;
        RECT 150.480 8.380 150.830 10.540 ;
        RECT 154.630 7.900 154.800 63.420 ;
        RECT 149.830 7.730 154.800 7.900 ;
      LAYER mcon ;
        RECT 152.060 222.330 152.350 222.500 ;
        RECT 151.750 220.655 151.920 222.035 ;
        RECT 152.490 220.655 152.660 222.035 ;
        RECT 152.060 220.190 152.350 220.360 ;
        RECT 156.060 222.330 156.350 222.500 ;
        RECT 155.750 220.655 155.920 222.035 ;
        RECT 156.490 220.655 156.660 222.035 ;
        RECT 156.060 220.190 156.350 220.360 ;
        RECT 152.060 218.240 152.350 218.410 ;
        RECT 151.750 217.110 151.920 217.990 ;
        RECT 152.490 217.110 152.660 217.990 ;
        RECT 152.060 216.690 152.350 216.860 ;
        RECT 156.060 218.240 156.350 218.410 ;
        RECT 155.750 217.110 155.920 217.990 ;
        RECT 156.490 217.110 156.660 217.990 ;
        RECT 156.060 216.690 156.350 216.860 ;
        RECT 149.060 197.740 156.900 197.910 ;
        RECT 148.750 190.610 148.920 197.490 ;
        RECT 157.040 190.610 157.210 197.490 ;
        RECT 149.060 190.190 156.900 190.360 ;
        RECT 150.560 168.740 158.400 168.910 ;
        RECT 150.250 161.610 150.420 168.490 ;
        RECT 158.540 161.610 158.710 168.490 ;
        RECT 150.560 161.190 158.400 161.360 ;
        RECT 151.560 127.740 159.400 127.910 ;
        RECT 151.250 120.610 151.420 127.490 ;
        RECT 159.540 120.610 159.710 127.490 ;
        RECT 151.560 120.190 159.400 120.360 ;
        RECT 151.060 86.240 158.900 86.410 ;
        RECT 150.750 79.110 150.920 85.990 ;
        RECT 159.040 79.110 159.210 85.990 ;
        RECT 151.060 78.690 158.900 78.860 ;
      LAYER met1 ;
        RECT 152.000 222.300 152.410 222.530 ;
        RECT 156.000 222.300 156.410 222.530 ;
        RECT 151.720 220.595 151.950 222.095 ;
        RECT 152.460 220.595 152.690 222.095 ;
        RECT 155.720 220.595 155.950 222.095 ;
        RECT 156.460 220.595 156.690 222.095 ;
        RECT 152.000 220.160 152.410 220.390 ;
        RECT 156.000 220.160 156.410 220.390 ;
        RECT 152.000 218.210 152.410 218.440 ;
        RECT 156.000 218.210 156.410 218.440 ;
        RECT 151.720 217.050 151.950 218.050 ;
        RECT 152.460 217.050 152.690 218.050 ;
        RECT 155.720 217.050 155.950 218.050 ;
        RECT 156.460 217.050 156.690 218.050 ;
        RECT 152.000 216.660 152.410 216.890 ;
        RECT 156.000 216.660 156.410 216.890 ;
        RECT 149.000 197.710 156.960 197.940 ;
        RECT 148.720 190.550 148.950 197.550 ;
        RECT 157.010 190.550 157.240 197.550 ;
        RECT 149.000 190.160 156.960 190.390 ;
        RECT 150.500 168.710 158.460 168.940 ;
        RECT 150.220 161.550 150.450 168.550 ;
        RECT 158.510 161.550 158.740 168.550 ;
        RECT 150.500 161.160 158.460 161.390 ;
        RECT 151.500 127.710 159.460 127.940 ;
        RECT 151.220 120.550 151.450 127.550 ;
        RECT 159.510 120.550 159.740 127.550 ;
        RECT 151.500 120.160 159.460 120.390 ;
        RECT 151.000 86.210 158.960 86.440 ;
        RECT 150.720 79.050 150.950 86.050 ;
        RECT 159.010 79.050 159.240 86.050 ;
        RECT 151.000 78.660 158.960 78.890 ;
        RECT 148.020 8.780 148.430 8.840 ;
        RECT 150.450 8.780 150.860 8.840 ;
        RECT 148.020 8.380 150.860 8.780 ;
        RECT 148.020 8.320 148.430 8.380 ;
        RECT 150.450 8.320 150.860 8.380 ;
      LAYER via ;
        RECT 148.860 8.390 149.460 8.760 ;
      LAYER met2 ;
        RECT 148.860 8.340 149.460 8.810 ;
      LAYER via2 ;
        RECT 148.860 8.390 149.460 8.760 ;
      LAYER met3 ;
        RECT 109.500 187.000 135.995 213.000 ;
        RECT 104.000 153.500 130.495 179.500 ;
        RECT 104.000 115.000 130.495 141.000 ;
        RECT 99.500 76.500 130.995 102.500 ;
        RECT 148.810 8.365 149.510 8.785 ;
      LAYER via3 ;
        RECT 135.575 187.140 135.895 212.860 ;
        RECT 130.075 153.640 130.395 179.360 ;
        RECT 130.075 115.140 130.395 140.860 ;
        RECT 130.575 76.640 130.895 102.360 ;
        RECT 148.860 8.390 149.460 8.760 ;
      LAYER met4 ;
        RECT 4.290 224.760 4.295 225.760 ;
        RECT 3.995 224.005 4.295 224.760 ;
        RECT 7.670 224.005 7.970 224.760 ;
        RECT 11.350 224.005 11.650 224.760 ;
        RECT 15.030 224.005 15.330 224.760 ;
        RECT 18.710 224.005 19.010 224.760 ;
        RECT 22.390 224.005 22.690 224.760 ;
        RECT 26.070 224.005 26.370 224.760 ;
        RECT 29.750 224.005 30.050 224.760 ;
        RECT 33.430 224.005 33.730 224.760 ;
        RECT 37.110 224.005 37.410 224.760 ;
        RECT 40.790 224.005 41.090 224.760 ;
        RECT 44.470 224.005 44.770 224.760 ;
        RECT 48.150 224.005 48.450 224.760 ;
        RECT 51.830 224.005 52.130 224.760 ;
        RECT 55.510 224.005 55.810 224.760 ;
        RECT 59.190 224.005 59.490 224.760 ;
        RECT 62.870 224.005 63.170 224.760 ;
        RECT 66.550 224.005 66.850 224.760 ;
        RECT 70.230 224.005 70.530 224.760 ;
        RECT 73.910 224.005 74.210 224.760 ;
        RECT 77.590 224.005 77.890 224.760 ;
        RECT 81.270 224.005 81.570 224.760 ;
        RECT 84.950 224.005 85.250 224.760 ;
        RECT 88.630 224.005 88.930 224.760 ;
        RECT 3.995 223.705 88.945 224.005 ;
        RECT 49.000 220.760 50.500 223.705 ;
        RECT 84.950 223.700 85.250 223.705 ;
        RECT 88.630 223.700 88.930 223.705 ;
        RECT 110.195 187.695 134.805 212.305 ;
        RECT 135.495 187.060 135.975 212.940 ;
        RECT 104.695 154.195 129.305 178.805 ;
        RECT 129.995 153.560 130.475 179.440 ;
        RECT 104.695 115.695 129.305 140.305 ;
        RECT 129.995 115.060 130.475 140.940 ;
        RECT 100.195 77.195 129.805 101.805 ;
        RECT 130.495 76.560 130.975 102.440 ;
        RECT 148.850 8.765 149.450 8.790 ;
        RECT 148.850 8.385 149.465 8.765 ;
        RECT 148.850 7.250 149.450 8.385 ;
        RECT 148.850 6.650 157.160 7.250 ;
        RECT 156.560 1.000 157.160 6.650 ;
  END
END tt_um_urish_charge_pump
END LIBRARY

