magic
tech sky130A
magscale 1 2
timestamp 1711889643
<< error_s >>
rect 19900 43054 22280 43340
rect 19900 41366 20186 43054
rect 21994 41366 22280 43054
rect 19900 41080 22280 41366
rect 19840 37474 22220 37760
rect 19840 35786 20126 37474
rect 21934 35786 22220 37474
rect 19840 35500 22220 35786
rect 19840 32014 22220 32300
rect 19840 30326 20126 32014
rect 21934 30326 22220 32014
rect 19840 30040 22220 30326
<< dnwell >>
rect 19980 41160 22200 43260
rect 19920 35580 22140 37680
rect 19920 30120 22140 32220
<< locali >>
rect 31012 43728 31070 43762
<< viali >>
rect 30512 44468 30570 44502
rect 31012 44466 31070 44500
rect 31212 44302 31246 44356
rect 31212 43542 31246 43596
rect 21542 43050 21602 43084
rect 20160 37440 20340 37500
rect 20160 31980 20340 32040
rect 29610 1676 29680 1756
rect 30096 1676 30166 1756
<< metal1 >>
rect 30500 44502 30760 44520
rect 30500 44468 30512 44502
rect 30570 44468 30760 44502
rect 30500 44460 30760 44468
rect 30820 44506 31080 44520
rect 30820 44500 31082 44506
rect 30820 44466 31012 44500
rect 31070 44466 31082 44500
rect 30820 44460 31082 44466
rect 31200 44360 31260 44520
rect 29150 44280 29160 44340
rect 29340 44280 30480 44340
rect 30580 44300 31000 44360
rect 31100 44356 31260 44360
rect 31100 44302 31212 44356
rect 31246 44302 31260 44356
rect 31100 44300 31260 44302
rect 30760 43980 30820 44300
rect 30750 43920 30760 43980
rect 30820 43920 30830 43980
rect 30760 43780 30820 43920
rect 30480 43720 31100 43780
rect 29150 43620 29160 43680
rect 29340 43620 30480 43680
rect 31200 43600 31260 44300
rect 30600 43540 30980 43600
rect 31100 43596 31260 43600
rect 31100 43542 31212 43596
rect 31246 43542 31260 43596
rect 31100 43540 31260 43542
rect 21470 43260 21480 43440
rect 21660 43260 21670 43440
rect 21480 43090 21600 43260
rect 21480 43084 21614 43090
rect 21480 43050 21542 43084
rect 21602 43050 21614 43084
rect 21480 43044 21614 43050
rect 21480 43020 21600 43044
rect 20220 42960 21600 43020
rect 30680 42960 30740 43540
rect 31200 43400 31260 43540
rect 31190 43280 31200 43400
rect 31260 43280 31270 43400
rect 20220 42900 20340 42960
rect 20220 42720 20280 42900
rect 21900 42120 22140 42300
rect 22320 42120 22330 42300
rect 20150 37680 20160 37860
rect 20340 37680 20350 37860
rect 20160 37506 20340 37680
rect 20148 37500 20352 37506
rect 20148 37440 20160 37500
rect 20340 37440 20352 37500
rect 20148 37434 20352 37440
rect 20160 37140 20340 37434
rect 21840 36480 22140 36660
rect 22320 36480 22330 36660
rect 20150 32220 20160 32400
rect 20340 32220 20350 32400
rect 20160 32046 20340 32220
rect 20148 32040 20352 32046
rect 20148 31980 20160 32040
rect 20340 31980 20352 32040
rect 20148 31974 20352 31980
rect 20160 31680 20340 31974
rect 21840 31080 22140 31260
rect 22320 31080 22330 31260
rect 29604 1756 29686 1768
rect 30090 1756 30172 1768
rect 29604 1676 29610 1756
rect 29680 1752 30096 1756
rect 29680 1678 29772 1752
rect 29892 1678 30096 1752
rect 29680 1676 30096 1678
rect 30166 1676 30172 1756
rect 29604 1664 29686 1676
rect 30090 1664 30172 1676
<< via1 >>
rect 30760 44460 30820 44520
rect 29160 44280 29340 44340
rect 30760 43920 30820 43980
rect 29160 43620 29340 43680
rect 21480 43260 21660 43440
rect 31200 43280 31260 43400
rect 22140 42120 22320 42300
rect 20160 37680 20340 37860
rect 22140 36480 22320 36660
rect 20160 32220 20340 32400
rect 22140 31080 22320 31260
rect 29772 1678 29892 1752
<< metal2 >>
rect 30760 44940 30820 44950
rect 30760 44520 30820 44860
rect 30760 44450 30820 44460
rect 29160 44340 29340 44350
rect 29160 44270 29340 44280
rect 27900 43980 28020 43990
rect 30760 43980 30820 43990
rect 28020 43920 30760 43980
rect 30820 43920 30840 43980
rect 28020 43860 30840 43920
rect 27900 43850 28020 43860
rect 29160 43680 29340 43690
rect 29160 43610 29340 43620
rect 21480 43440 21660 43450
rect 31200 43400 31260 43410
rect 31200 43270 31260 43280
rect 21480 43250 21660 43260
rect 22140 42300 22320 42310
rect 20160 37860 20340 37870
rect 22140 37860 22320 42120
rect 20340 37680 22320 37860
rect 20160 37670 20340 37680
rect 22140 36660 22320 36670
rect 20160 32400 20340 32410
rect 22140 32400 22320 36480
rect 20340 32220 22320 32400
rect 20160 32210 20340 32220
rect 22140 31260 22320 31270
rect 22140 31070 22320 31080
rect 29772 1752 29892 1762
rect 29772 1668 29892 1678
<< via2 >>
rect 30760 44860 30820 44940
rect 29160 44280 29340 44340
rect 27900 43860 28020 43980
rect 29160 43620 29340 43680
rect 21480 43260 21660 43440
rect 31200 43280 31260 43400
rect 22140 42120 22320 42300
rect 22140 36480 22320 36660
rect 22140 31080 22320 31260
rect 29772 1678 29892 1752
<< metal3 >>
rect 30750 44940 30830 44945
rect 30730 44860 30740 44940
rect 30840 44860 30850 44940
rect 30750 44855 30830 44860
rect 29090 44500 29100 44800
rect 29400 44500 29410 44800
rect 29100 44340 29400 44500
rect 29100 44280 29160 44340
rect 29340 44280 29400 44340
rect 27890 43980 28030 43985
rect 27890 43860 27900 43980
rect 28020 43860 28030 43980
rect 27890 43855 28030 43860
rect 29100 43680 29400 44280
rect 29100 43620 29160 43680
rect 29340 43620 29400 43680
rect 29100 43600 29400 43620
rect 21470 43440 21670 43445
rect 21420 43260 21480 43440
rect 21660 43260 28200 43440
rect 28500 43400 28510 43440
rect 31190 43400 31270 43405
rect 28500 43280 31200 43400
rect 31260 43280 31270 43400
rect 28500 43260 28510 43280
rect 31190 43275 31270 43280
rect 21470 43255 21670 43260
rect 22130 42300 22330 42305
rect 22130 42120 22140 42300
rect 22320 42120 22330 42300
rect 22130 42115 22330 42120
rect 22130 36660 22330 36665
rect 22130 36480 22140 36660
rect 22320 36480 22330 36660
rect 22130 36475 22330 36480
rect 22130 31260 22330 31265
rect 22130 31080 22140 31260
rect 22320 31080 22330 31260
rect 22130 31075 22330 31080
rect 29762 1752 29902 1757
rect 29762 1678 29772 1752
rect 29892 1678 29902 1752
rect 29762 1673 29902 1678
<< via3 >>
rect 30740 44860 30760 44940
rect 30760 44860 30820 44940
rect 30820 44860 30840 44940
rect 29100 44500 29400 44800
rect 27900 43860 28020 43980
rect 28200 43260 28500 43440
rect 22140 42120 22320 42300
rect 22140 36480 22320 36660
rect 22140 31080 22320 31260
rect 29772 1678 29892 1752
<< metal4 >>
rect 798 44952 859 45152
rect 799 44801 859 44952
rect 1534 44801 1594 45152
rect 2270 44801 2330 45152
rect 3006 44801 3066 45152
rect 3742 44801 3802 45152
rect 4478 44801 4538 45152
rect 5214 44801 5274 45152
rect 5950 44801 6010 45152
rect 6686 44801 6746 45152
rect 7422 44801 7482 45152
rect 8158 44801 8218 45152
rect 8894 44801 8954 45152
rect 9630 44801 9690 45152
rect 10366 44801 10426 45152
rect 11102 44801 11162 45152
rect 11838 44801 11898 45152
rect 12574 44801 12634 45152
rect 13310 44801 13370 45152
rect 14046 44801 14106 45152
rect 14782 44801 14842 45152
rect 15518 44801 15578 45152
rect 16254 44801 16314 45152
rect 16990 44801 17050 45152
rect 17726 44801 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30739 44940 30841 44941
rect 30739 44860 30740 44940
rect 30840 44930 30841 44940
rect 30974 44930 31034 45152
rect 31710 44952 31770 45152
rect 30840 44870 31034 44930
rect 30840 44860 30841 44870
rect 30739 44859 30841 44860
rect 799 44800 17789 44801
rect 29099 44800 29401 44801
rect 799 44741 29100 44800
rect 800 44700 29100 44741
rect 9800 44500 29100 44700
rect 29400 44500 29401 44800
rect 9800 27840 10100 44500
rect 29099 44499 29401 44500
rect 27899 43980 28021 43981
rect 27899 43860 27900 43980
rect 28020 43860 28021 43980
rect 27899 43859 28021 43860
rect 27900 43020 28020 43859
rect 28200 43441 28500 44152
rect 28199 43440 28501 43441
rect 28199 43260 28200 43440
rect 28500 43260 28501 43440
rect 28199 43259 28501 43260
rect 22139 42300 22321 42301
rect 22139 42120 22140 42300
rect 22320 42120 22920 42300
rect 22139 42119 22321 42120
rect 22139 36660 22321 36661
rect 22139 36480 22140 36660
rect 22320 36480 22860 36660
rect 22139 36479 22321 36480
rect 22139 31260 22321 31261
rect 22139 31080 22140 31260
rect 22320 31080 22860 31260
rect 22139 31079 22321 31080
rect 9800 25680 13560 27840
rect 9800 1000 10100 25680
rect 28200 1000 28500 43259
rect 29770 1753 29890 1758
rect 29770 1752 29893 1753
rect 29770 1678 29772 1752
rect 29892 1678 29893 1752
rect 29770 1677 29893 1678
rect 29770 1450 29890 1677
rect 29770 1330 31432 1450
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 1330
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C1
timestamp 1711870259
transform 1 0 25350 0 1 40500
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C2
timestamp 1711870259
transform 1 0 25330 0 1 35060
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C3
timestamp 1711870259
transform 1 0 25330 0 1 29600
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_WMZ6NR  C4
timestamp 1711870259
transform 1 0 16410 0 1 26600
box -3150 -2600 3149 2600
use sky130_fd_pr__pfet_01v8_BFP3TE  M1
timestamp 1711870259
transform 1 0 31041 0 1 44269
box -241 -369 241 369
use sky130_fd_pr__pfet_01v8_BFP3TE  M2
timestamp 1711870259
transform 1 0 31041 0 1 43531
box -241 -369 241 369
use sky130_fd_pr__nfet_01v8_DSY3K9  M3
timestamp 1711870259
transform -1 0 30541 0 1 44330
box -241 -310 241 310
use sky130_fd_pr__nfet_01v8_DSY3K9  M4
timestamp 1711870259
transform 1 0 30541 0 1 43592
box -241 -310 241 310
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M5
timestamp 1711870259
transform 1 0 21096 0 1 42210
box -996 -910 996 910
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M6
timestamp 1711870259
transform 1 0 21036 0 1 36610
box -996 -910 996 910
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M7
timestamp 1711870259
transform 1 0 21036 0 1 31150
box -996 -910 996 910
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M8
timestamp 1711870259
transform 1 0 21036 0 1 28330
box -996 -910 996 910
use sky130_fd_pr__res_xhigh_po_0p35_5JC923  R1
timestamp 1711870259
transform 1 0 30463 0 1 7132
box -533 -5622 533 5622
use sky130_fd_pr__res_xhigh_po_0p35_VR8WVB  R2
timestamp 1711870259
transform 1 0 25578 0 1 6846
box -4268 -5336 4268 5336
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 28200 1000 28500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 30760 43980 30820 44100 0 FreeSans 320 90 0 0 clka
flabel metal1 30680 42960 30740 43560 0 FreeSans 320 90 0 0 clkb
flabel metal2 22140 37800 22320 42120 0 FreeSans 1600 0 0 0 stage1
flabel metal2 22140 32400 22320 36480 0 FreeSans 1600 0 0 0 stage2
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
