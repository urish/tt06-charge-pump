magic
tech sky130A
magscale 1 2
timestamp 1711870259
<< metal3 >>
rect -2650 2572 2649 2600
rect -2650 -2572 2565 2572
rect 2629 -2572 2649 2572
rect -2650 -2600 2649 -2572
<< via3 >>
rect 2565 -2572 2629 2572
<< mimcap >>
rect -2550 2460 2450 2500
rect -2550 -2460 -2510 2460
rect 2410 -2460 2450 2460
rect -2550 -2500 2450 -2460
<< mimcapcontact >>
rect -2510 -2460 2410 2460
<< metal4 >>
rect 2549 2572 2645 2588
rect -2511 2460 2411 2461
rect -2511 -2460 -2510 2460
rect 2410 -2460 2411 2460
rect -2511 -2461 2411 -2460
rect 2549 -2572 2565 2572
rect 2629 -2572 2645 2572
rect 2549 -2588 2645 -2572
<< properties >>
string FIXED_BBOX -2650 -2600 2550 2600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
