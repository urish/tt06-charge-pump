magic
tech sky130A
magscale 1 2
timestamp 1711870259
<< pwell >>
rect -533 -5622 533 5622
<< psubdiff >>
rect -497 5552 -401 5586
rect 401 5552 497 5586
rect -497 5490 -463 5552
rect 463 5490 497 5552
rect -497 -5552 -463 -5490
rect 463 -5552 497 -5490
rect -497 -5586 -401 -5552
rect 401 -5586 497 -5552
<< psubdiffcont >>
rect -401 5552 401 5586
rect -497 -5490 -463 5490
rect 463 -5490 497 5490
rect -401 -5586 401 -5552
<< xpolycontact >>
rect 297 5024 367 5456
rect -367 -5456 -297 -5024
<< xpolyres >>
rect -367 4850 -131 4920
rect -367 -5024 -297 4850
rect -201 -4850 -131 4850
rect -35 4850 201 4920
rect -35 -4850 35 4850
rect -201 -4920 35 -4850
rect 131 -4850 201 4850
rect 297 -4850 367 5024
rect 131 -4920 367 -4850
<< locali >>
rect -497 5552 -401 5586
rect 401 5552 497 5586
rect -497 5490 -463 5552
rect 463 5490 497 5552
rect -497 -5552 -463 -5490
rect 463 -5552 497 -5490
rect -497 -5586 -401 -5552
rect 401 -5586 497 -5552
<< properties >>
string FIXED_BBOX -480 -5569 480 5569
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 49.2 m 1 nx 5 wmin 0.350 lmin 0.50 rho 2000 val 1.414meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
