magic
tech sky130A
timestamp 1711967973
<< metal2 >>
rect 1540 2856 1736 2884
rect 1512 2828 1764 2856
rect 1512 2800 1792 2828
rect 1484 2772 1792 2800
rect 1484 2744 1820 2772
rect 1456 2716 1820 2744
rect 1428 2688 1848 2716
rect 1428 2660 1876 2688
rect 1400 2632 1876 2660
rect 1400 2604 1904 2632
rect 1372 2576 1904 2604
rect 1372 2548 1932 2576
rect 1344 2520 1932 2548
rect 5880 2520 5992 2548
rect 1316 2492 1960 2520
rect 5796 2492 6076 2520
rect 1316 2464 1988 2492
rect 5768 2464 6104 2492
rect 1288 2436 1988 2464
rect 1288 2408 1624 2436
rect 1652 2408 2016 2436
rect 5740 2408 6132 2464
rect 1260 2380 1624 2408
rect 1680 2380 2016 2408
rect 1260 2352 1596 2380
rect 1680 2352 2044 2380
rect 1232 2324 1568 2352
rect 1708 2324 2044 2352
rect 1204 2296 1568 2324
rect 1736 2296 2072 2324
rect 1204 2268 1540 2296
rect 1736 2268 2100 2296
rect 1176 2240 1540 2268
rect 1764 2240 2100 2268
rect 1176 2212 1512 2240
rect 1764 2212 2128 2240
rect 1148 2184 1484 2212
rect 1120 2156 1484 2184
rect 1792 2184 2128 2212
rect 1792 2156 2156 2184
rect 1120 2128 1456 2156
rect 1820 2128 2156 2156
rect 1092 2100 1456 2128
rect 1848 2100 2184 2128
rect 1092 2072 1428 2100
rect 1848 2072 2212 2100
rect 1064 2044 1428 2072
rect 1876 2044 2212 2072
rect 1064 2016 1400 2044
rect 1876 2016 2240 2044
rect 1036 1988 1372 2016
rect 1904 1988 2240 2016
rect 1008 1960 1372 1988
rect 1008 1932 1344 1960
rect 980 1904 1344 1932
rect 1484 1904 1820 1988
rect 1932 1960 2268 1988
rect 1932 1932 2296 1960
rect 1960 1904 2296 1932
rect 980 1876 1316 1904
rect 1484 1876 1792 1904
rect 1960 1876 2324 1904
rect 952 1848 1316 1876
rect 1456 1848 1792 1876
rect 1988 1848 2324 1876
rect 952 1820 1288 1848
rect 924 1792 1260 1820
rect 1456 1792 1764 1848
rect 1988 1820 2352 1848
rect 2016 1792 2352 1820
rect 896 1764 1260 1792
rect 1428 1764 1764 1792
rect 2044 1764 2380 1792
rect 896 1736 1232 1764
rect 868 1708 1232 1736
rect 1428 1708 1736 1764
rect 2044 1736 2408 1764
rect 2072 1708 2408 1736
rect 868 1680 1204 1708
rect 1428 1680 1708 1708
rect 2072 1680 2436 1708
rect 840 1652 1204 1680
rect 840 1624 1176 1652
rect 1400 1624 1708 1680
rect 2100 1652 2436 1680
rect 3836 1652 4172 2352
rect 4732 1652 5068 2352
rect 5712 2240 6160 2408
rect 5740 2184 6132 2240
rect 5768 2156 6104 2184
rect 5796 2128 6076 2156
rect 5852 2100 6020 2128
rect 7168 1960 7560 1988
rect 5404 1708 6132 1960
rect 7084 1932 8036 1960
rect 7028 1904 8036 1932
rect 7000 1876 8036 1904
rect 6944 1848 8036 1876
rect 6916 1792 8036 1848
rect 6888 1764 8036 1792
rect 6860 1736 8036 1764
rect 6860 1708 7252 1736
rect 7476 1708 8036 1736
rect 8288 1848 8624 2492
rect 11032 2296 11424 2352
rect 12152 2296 12516 2352
rect 11032 2268 11452 2296
rect 11060 2184 11452 2268
rect 12124 2240 12516 2296
rect 12124 2184 12488 2240
rect 14196 2212 14924 2492
rect 16072 2352 16212 2380
rect 15988 2324 16212 2352
rect 15876 2296 16212 2324
rect 11088 2100 11480 2184
rect 12096 2156 12488 2184
rect 12096 2100 12460 2156
rect 11116 1988 11508 2100
rect 12068 2072 12460 2100
rect 12068 1988 12432 2072
rect 8820 1960 9156 1988
rect 8764 1932 9212 1960
rect 8708 1904 9268 1932
rect 11144 1904 11536 1988
rect 8680 1876 9296 1904
rect 8652 1848 9324 1876
rect 8288 1792 9352 1848
rect 11172 1820 11564 1904
rect 12040 1876 12404 1988
rect 13048 1960 13468 1988
rect 12964 1932 13552 1960
rect 12908 1904 13608 1932
rect 12852 1876 13664 1904
rect 11200 1792 11564 1820
rect 12012 1792 12376 1876
rect 12824 1848 13692 1876
rect 12796 1820 13720 1848
rect 12768 1792 13748 1820
rect 8288 1708 9380 1792
rect 11200 1736 11592 1792
rect 2100 1624 2464 1652
rect 812 1596 1148 1624
rect 1400 1596 1680 1624
rect 2128 1596 2464 1624
rect 784 1568 1148 1596
rect 784 1540 1120 1568
rect 756 1512 1120 1540
rect 1372 1540 1680 1596
rect 2156 1568 2492 1596
rect 2156 1540 2520 1568
rect 756 1484 1092 1512
rect 1372 1484 1652 1540
rect 2184 1512 2520 1540
rect 2184 1484 2548 1512
rect 728 1456 1064 1484
rect 700 1428 1064 1456
rect 700 1400 1036 1428
rect 672 1372 1036 1400
rect 1344 1400 1624 1484
rect 1904 1456 1960 1484
rect 1848 1428 1960 1456
rect 2212 1456 2548 1484
rect 2212 1428 2576 1456
rect 1792 1400 1932 1428
rect 2240 1400 2576 1428
rect 1344 1372 1596 1400
rect 1736 1372 1932 1400
rect 672 1344 1008 1372
rect 644 1316 1008 1344
rect 1316 1316 1596 1372
rect 1680 1344 1932 1372
rect 2268 1372 2604 1400
rect 3836 1372 5068 1652
rect 2268 1344 2632 1372
rect 1624 1316 1904 1344
rect 644 1288 980 1316
rect 1316 1288 1904 1316
rect 2296 1316 2632 1344
rect 2296 1288 2660 1316
rect 616 1260 952 1288
rect 588 1232 952 1260
rect 1288 1232 1904 1288
rect 2324 1260 2660 1288
rect 2352 1232 2688 1260
rect 588 1204 924 1232
rect 560 1176 924 1204
rect 1288 1176 1876 1232
rect 2352 1204 2716 1232
rect 560 1148 896 1176
rect 532 1120 896 1148
rect 1260 1148 1624 1176
rect 1260 1120 1540 1148
rect 1652 1120 1876 1176
rect 2380 1176 2716 1204
rect 2380 1148 2744 1176
rect 2408 1120 2744 1148
rect 532 1092 868 1120
rect 1260 1092 1484 1120
rect 1652 1092 1848 1120
rect 2408 1092 2772 1120
rect 504 1064 840 1092
rect 1260 1064 1428 1092
rect 476 1036 840 1064
rect 1232 1036 1372 1064
rect 1624 1036 1848 1092
rect 2436 1064 2772 1092
rect 2464 1036 2800 1064
rect 476 1008 812 1036
rect 1232 1008 1316 1036
rect 448 980 812 1008
rect 448 952 784 980
rect 1624 952 1820 1036
rect 2464 1008 2828 1036
rect 2492 980 2828 1008
rect 2492 952 2856 980
rect 420 924 784 952
rect 1596 924 1820 952
rect 2520 924 2856 952
rect 420 896 756 924
rect 392 868 728 896
rect 364 840 728 868
rect 1596 840 1792 924
rect 2520 896 2884 924
rect 2548 868 2884 896
rect 2576 840 2912 868
rect 364 812 700 840
rect 336 784 700 812
rect 1596 784 1764 840
rect 2576 812 2940 840
rect 336 756 672 784
rect 1456 756 1512 784
rect 308 728 644 756
rect 1456 728 1540 756
rect 1568 728 1764 784
rect 2604 784 2940 812
rect 2604 756 2968 784
rect 2632 728 2968 756
rect 280 700 644 728
rect 280 672 616 700
rect 252 644 616 672
rect 1484 672 1736 728
rect 1820 700 1848 728
rect 2632 700 2996 728
rect 1764 672 1848 700
rect 2660 672 2996 700
rect 252 616 588 644
rect 1484 616 1820 672
rect 2688 644 3024 672
rect 2688 616 3052 644
rect 3836 616 4172 1372
rect 4732 616 5068 1372
rect 5768 896 6132 1708
rect 6832 1680 7224 1708
rect 7504 1680 7868 1708
rect 6832 1652 7196 1680
rect 7532 1652 7868 1680
rect 8288 1680 8904 1708
rect 8960 1680 9408 1708
rect 8288 1652 8820 1680
rect 9016 1652 9408 1680
rect 6832 1596 7168 1652
rect 6832 1456 7140 1596
rect 7560 1568 7896 1652
rect 7588 1484 7896 1568
rect 6832 1400 7168 1456
rect 7560 1400 7896 1484
rect 6832 1344 7196 1400
rect 7532 1372 7896 1400
rect 8288 1624 8792 1652
rect 8288 1596 8764 1624
rect 9044 1596 9408 1652
rect 11228 1680 11592 1736
rect 11984 1708 12348 1792
rect 12740 1764 13776 1792
rect 12712 1736 13776 1764
rect 12712 1708 13804 1736
rect 11984 1680 12320 1708
rect 12684 1680 13216 1708
rect 13272 1680 13804 1708
rect 11228 1624 11620 1680
rect 8288 1568 8736 1596
rect 8288 1540 8708 1568
rect 8288 1512 8680 1540
rect 8288 1484 8652 1512
rect 7504 1344 7868 1372
rect 6860 1316 7252 1344
rect 7476 1316 7868 1344
rect 6860 1288 7868 1316
rect 6888 1260 7840 1288
rect 6916 1232 7812 1260
rect 6916 1204 7784 1232
rect 6888 1176 7756 1204
rect 6860 1148 7728 1176
rect 6860 1120 7700 1148
rect 6832 1092 7644 1120
rect 6832 1064 7140 1092
rect 7196 1064 7532 1092
rect 6804 952 7112 1064
rect 6804 924 7168 952
rect 6804 896 7224 924
rect 5348 616 6524 896
rect 6804 868 7700 896
rect 6804 840 7784 868
rect 6832 812 7868 840
rect 6832 784 7896 812
rect 6860 756 7952 784
rect 6888 700 7980 756
rect 6860 672 8008 700
rect 6832 644 8008 672
rect 6804 616 7196 644
rect 7476 616 8036 644
rect 8288 616 8624 1484
rect 9072 616 9408 1596
rect 11256 1596 11620 1624
rect 11956 1624 12320 1680
rect 12656 1652 13132 1680
rect 13384 1652 13832 1680
rect 12656 1624 13076 1652
rect 13412 1624 13832 1652
rect 11956 1596 12292 1624
rect 12656 1596 13048 1624
rect 13440 1596 13860 1624
rect 11256 1540 11648 1596
rect 11284 1484 11648 1540
rect 11928 1512 12292 1596
rect 12628 1540 13020 1596
rect 13468 1568 13860 1596
rect 13496 1540 13860 1568
rect 12628 1512 12992 1540
rect 11928 1484 12264 1512
rect 11284 1456 11676 1484
rect 11312 1400 11676 1456
rect 11900 1428 12264 1484
rect 12600 1484 12992 1512
rect 13496 1484 13888 1540
rect 11900 1400 12236 1428
rect 11312 1344 11704 1400
rect 11340 1288 11704 1344
rect 11872 1344 12236 1400
rect 11872 1288 12208 1344
rect 11340 1260 11732 1288
rect 11368 1176 11732 1260
rect 11844 1260 12208 1288
rect 12600 1316 12964 1484
rect 12600 1260 12936 1316
rect 11844 1204 12180 1260
rect 11396 1092 11760 1176
rect 11816 1148 12180 1204
rect 11816 1092 12152 1148
rect 11424 1064 12152 1092
rect 12600 1092 12964 1260
rect 13524 1120 13888 1484
rect 13496 1092 13888 1120
rect 11424 980 12124 1064
rect 12600 1036 12992 1092
rect 13496 1036 13860 1092
rect 12628 980 13020 1036
rect 13468 1008 13860 1036
rect 13440 980 13860 1008
rect 11452 896 12096 980
rect 12628 952 13048 980
rect 13440 952 13832 980
rect 12656 924 13104 952
rect 13384 924 13832 952
rect 12656 896 13160 924
rect 13356 896 13804 924
rect 14560 896 14924 2212
rect 15848 1960 16212 2296
rect 17360 1960 17864 1988
rect 18900 1960 19292 1988
rect 20412 1960 20804 1988
rect 15512 1708 16716 1960
rect 17248 1932 17976 1960
rect 18816 1932 19768 1960
rect 20328 1932 20860 1960
rect 17164 1904 18032 1932
rect 18760 1904 19768 1932
rect 20272 1904 20916 1932
rect 17136 1876 18060 1904
rect 18704 1876 19768 1904
rect 20216 1876 20972 1904
rect 17136 1848 18088 1876
rect 18676 1848 19768 1876
rect 20188 1848 21000 1876
rect 17136 1820 18116 1848
rect 18648 1820 19768 1848
rect 20160 1820 21028 1848
rect 17136 1764 18144 1820
rect 18620 1764 19768 1820
rect 20132 1792 21056 1820
rect 20104 1764 21084 1792
rect 17136 1736 18172 1764
rect 18592 1736 19768 1764
rect 17136 1708 17472 1736
rect 17696 1708 18172 1736
rect 15848 1008 16212 1708
rect 17136 1680 17332 1708
rect 17752 1680 18172 1708
rect 18564 1708 18984 1736
rect 19180 1708 19768 1736
rect 20076 1736 21084 1764
rect 20076 1708 20524 1736
rect 20664 1708 21112 1736
rect 18564 1680 18928 1708
rect 19236 1680 19572 1708
rect 20048 1680 20440 1708
rect 20720 1680 21112 1708
rect 17136 1652 17248 1680
rect 17808 1652 18200 1680
rect 17136 1624 17192 1652
rect 17836 1568 18200 1652
rect 18564 1624 18900 1680
rect 19264 1624 19600 1680
rect 20048 1652 20412 1680
rect 20748 1652 21140 1680
rect 20020 1624 20384 1652
rect 20776 1624 21140 1652
rect 17864 1456 18200 1568
rect 17472 1428 18200 1456
rect 17360 1400 18200 1428
rect 18536 1428 18872 1624
rect 19292 1428 19628 1624
rect 20020 1596 20356 1624
rect 19992 1568 20356 1596
rect 19992 1484 20328 1568
rect 20804 1540 21168 1624
rect 19964 1456 20328 1484
rect 20832 1456 21168 1540
rect 18536 1400 18900 1428
rect 17276 1372 18200 1400
rect 17220 1344 18200 1372
rect 17192 1316 18200 1344
rect 18564 1372 18900 1400
rect 19264 1372 19600 1428
rect 18564 1344 18928 1372
rect 19236 1344 19600 1372
rect 18564 1316 18984 1344
rect 19180 1316 19600 1344
rect 17164 1288 18200 1316
rect 18592 1288 19572 1316
rect 17136 1260 18200 1288
rect 17108 1232 18200 1260
rect 17080 1204 18200 1232
rect 17080 1176 17556 1204
rect 17052 1148 17500 1176
rect 17052 1120 17444 1148
rect 17052 1092 17416 1120
rect 17024 1064 17416 1092
rect 15876 952 16240 1008
rect 17024 980 17388 1064
rect 17864 1036 18200 1204
rect 18620 1260 19572 1288
rect 18620 1232 19544 1260
rect 18620 1204 19516 1232
rect 19964 1204 21168 1456
rect 18620 1176 19488 1204
rect 18592 1148 19460 1176
rect 18564 1120 19404 1148
rect 19964 1120 20300 1204
rect 18564 1092 19348 1120
rect 17836 1008 18200 1036
rect 18536 1064 18872 1092
rect 18928 1064 19264 1092
rect 19964 1064 20328 1120
rect 18536 1036 18844 1064
rect 19964 1036 20356 1064
rect 18536 1008 18816 1036
rect 19992 1008 20356 1036
rect 17808 980 18200 1008
rect 17024 952 17416 980
rect 17752 952 18200 980
rect 15876 924 16268 952
rect 17052 924 17416 952
rect 17724 924 18200 952
rect 15876 896 16296 924
rect 16688 896 16716 924
rect 11480 868 12096 896
rect 12684 868 13804 896
rect 11480 812 12068 868
rect 12684 840 13776 868
rect 11508 784 12068 812
rect 12712 784 13748 840
rect 11508 728 12040 784
rect 12740 756 13720 784
rect 12768 728 13692 756
rect 11536 700 12040 728
rect 12796 700 13636 728
rect 11536 616 12012 700
rect 12852 672 13608 700
rect 12908 644 13552 672
rect 12964 616 13496 644
rect 14140 616 15316 896
rect 15876 868 16352 896
rect 16548 868 16716 896
rect 15876 840 16716 868
rect 15904 784 16716 840
rect 17052 896 17444 924
rect 17696 896 18200 924
rect 17052 868 17500 896
rect 17640 868 18200 896
rect 18508 952 18844 1008
rect 19992 980 20384 1008
rect 19992 952 20412 980
rect 18508 924 18872 952
rect 20020 924 20440 952
rect 18508 896 18928 924
rect 20020 896 20496 924
rect 21000 896 21112 924
rect 18508 868 19404 896
rect 20048 868 20580 896
rect 20832 868 21112 896
rect 17052 812 18200 868
rect 18536 840 19516 868
rect 20048 840 21112 868
rect 18536 812 19572 840
rect 20076 812 21112 840
rect 15932 728 16716 784
rect 17080 756 18200 812
rect 18564 784 19628 812
rect 18564 756 19656 784
rect 20104 756 21112 812
rect 17108 728 17864 756
rect 15960 700 16716 728
rect 17136 700 17836 728
rect 15988 672 16716 700
rect 17164 672 17808 700
rect 16044 644 16716 672
rect 17192 644 17752 672
rect 16100 616 16716 644
rect 17248 616 17696 644
rect 17892 616 18200 756
rect 18592 728 19684 756
rect 20160 728 21112 756
rect 18620 700 19712 728
rect 20188 700 21112 728
rect 18592 672 19712 700
rect 20216 672 21112 700
rect 18536 644 19740 672
rect 20272 644 21112 672
rect 18536 616 18928 644
rect 19180 616 19740 644
rect 20328 616 21000 644
rect 224 588 588 616
rect 1512 588 1792 616
rect 2716 588 3052 616
rect 6776 588 7168 616
rect 7616 588 8036 616
rect 13076 588 13384 616
rect 16212 588 16548 616
rect 17332 588 17584 616
rect 18508 588 18900 616
rect 19320 588 19740 616
rect 20440 588 20832 616
rect 224 560 560 588
rect 196 532 532 560
rect 168 504 532 532
rect 1512 532 1764 588
rect 2716 560 3080 588
rect 6776 560 7140 588
rect 7644 560 8036 588
rect 2744 532 3080 560
rect 1512 504 1736 532
rect 2772 504 3108 532
rect 6748 504 7112 560
rect 168 476 504 504
rect 1512 476 1708 504
rect 2772 476 3136 504
rect 140 448 504 476
rect 1540 448 1708 476
rect 2800 448 3136 476
rect 140 420 476 448
rect 112 392 476 420
rect 1540 420 1680 448
rect 2800 420 3164 448
rect 112 364 448 392
rect 1540 364 1652 420
rect 2828 392 3164 420
rect 6748 420 7084 504
rect 7672 448 8036 560
rect 18480 532 18844 588
rect 19376 532 19768 588
rect 7644 420 8036 448
rect 6748 392 7112 420
rect 7644 392 8008 420
rect 2828 364 3192 392
rect 84 336 420 364
rect 1540 336 1624 364
rect 2856 336 3192 364
rect 6748 364 7140 392
rect 7616 364 8008 392
rect 6748 336 7196 364
rect 7532 336 8008 364
rect 18452 392 18816 532
rect 19404 476 19768 532
rect 19404 448 19740 476
rect 19376 420 19740 448
rect 19348 392 19740 420
rect 18452 364 18844 392
rect 19320 364 19740 392
rect 18452 336 18900 364
rect 19264 336 19712 364
rect 56 308 420 336
rect 1568 308 1596 336
rect 2884 308 3220 336
rect 6748 308 7336 336
rect 7392 308 7980 336
rect 18480 308 19040 336
rect 19124 308 19712 336
rect 56 280 392 308
rect 2884 280 3248 308
rect 28 252 3248 280
rect 6776 280 7952 308
rect 18480 280 19684 308
rect 6776 252 7924 280
rect 18508 252 19656 280
rect 28 224 3276 252
rect 6804 224 7896 252
rect 18508 224 19628 252
rect 0 196 3276 224
rect 6832 196 7868 224
rect 18536 196 19600 224
rect 0 84 3304 196
rect 6860 168 7840 196
rect 18592 168 19544 196
rect 6916 140 7784 168
rect 18620 140 19516 168
rect 6972 112 7728 140
rect 18704 112 19432 140
rect 7084 84 7616 112
rect 18788 84 19348 112
rect 0 56 3276 84
rect 28 28 3276 56
rect 28 0 3248 28
<< end >>
