VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_charge_pump
  CLASS BLOCK ;
  FOREIGN tt_um_urish_charge_pump ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.931599 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 142.200 5.000 143.700 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 151.500 220.100 153.910 223.200 ;
        RECT 151.500 216.410 153.910 219.510 ;
      LAYER nwell ;
        RECT 154.000 215.810 156.410 223.190 ;
        RECT 98.600 214.370 111.700 215.800 ;
        RECT 98.600 205.030 100.030 214.370 ;
      LAYER pwell ;
        RECT 100.200 205.200 110.160 214.300 ;
      LAYER nwell ;
        RECT 110.270 205.030 111.700 214.370 ;
        RECT 98.600 203.600 111.700 205.030 ;
        RECT 98.600 187.670 111.700 189.100 ;
        RECT 98.600 178.330 100.030 187.670 ;
      LAYER pwell ;
        RECT 100.200 178.500 110.160 187.600 ;
      LAYER nwell ;
        RECT 110.270 178.330 111.700 187.670 ;
        RECT 98.600 176.900 111.700 178.330 ;
        RECT 98.600 160.370 111.700 161.800 ;
        RECT 98.600 151.030 100.030 160.370 ;
      LAYER pwell ;
        RECT 100.200 151.200 110.160 160.300 ;
      LAYER nwell ;
        RECT 110.270 151.030 111.700 160.370 ;
        RECT 98.600 149.600 111.700 151.030 ;
        RECT 98.600 142.370 111.700 143.800 ;
        RECT 98.600 133.030 100.030 142.370 ;
      LAYER pwell ;
        RECT 100.200 133.200 110.160 142.300 ;
      LAYER nwell ;
        RECT 110.270 133.030 111.700 142.370 ;
        RECT 98.600 131.600 111.700 133.030 ;
      LAYER pwell ;
        RECT 106.550 7.550 149.230 60.910 ;
        RECT 149.650 7.550 159.130 60.990 ;
      LAYER li1 ;
        RECT 151.680 222.850 153.730 223.020 ;
        RECT 151.680 220.450 151.850 222.850 ;
        RECT 152.480 222.340 152.930 222.510 ;
        RECT 152.250 221.130 152.420 222.170 ;
        RECT 152.990 221.130 153.160 222.170 ;
        RECT 152.480 220.790 152.930 220.960 ;
        RECT 153.560 220.450 153.730 222.850 ;
        RECT 151.680 220.280 153.730 220.450 ;
        RECT 154.180 222.840 156.230 223.010 ;
        RECT 154.180 219.850 154.350 222.840 ;
        RECT 154.980 222.330 155.430 222.500 ;
        RECT 154.750 220.575 154.920 222.115 ;
        RECT 155.490 220.575 155.660 222.115 ;
        RECT 154.980 220.190 155.430 220.360 ;
        RECT 156.060 219.850 156.230 222.840 ;
        RECT 154.180 219.680 156.230 219.850 ;
        RECT 151.680 219.160 153.730 219.330 ;
        RECT 151.680 216.760 151.850 219.160 ;
        RECT 152.480 218.650 152.930 218.820 ;
        RECT 152.250 217.440 152.420 218.480 ;
        RECT 152.990 217.440 153.160 218.480 ;
        RECT 152.480 217.100 152.930 217.270 ;
        RECT 153.560 216.760 153.730 219.160 ;
        RECT 151.680 216.590 153.730 216.760 ;
        RECT 154.180 219.150 156.230 219.320 ;
        RECT 154.180 216.160 154.350 219.150 ;
        RECT 154.980 218.640 155.430 218.810 ;
        RECT 154.750 216.885 154.920 218.425 ;
        RECT 155.490 216.885 155.660 218.425 ;
        RECT 154.980 216.500 155.430 216.670 ;
        RECT 156.060 216.160 156.230 219.150 ;
        RECT 154.180 215.990 156.230 216.160 ;
        RECT 100.200 215.515 101.400 215.700 ;
        RECT 98.885 215.345 111.415 215.515 ;
        RECT 98.885 204.055 99.055 215.345 ;
        RECT 100.800 214.120 101.400 214.200 ;
        RECT 100.380 213.950 109.980 214.120 ;
        RECT 100.380 205.550 100.550 213.950 ;
        RECT 100.800 213.900 101.400 213.950 ;
        RECT 101.180 213.440 109.180 213.610 ;
        RECT 100.950 206.230 101.120 213.270 ;
        RECT 109.240 206.230 109.410 213.270 ;
        RECT 101.180 205.890 109.180 206.060 ;
        RECT 109.810 205.550 109.980 213.950 ;
        RECT 100.380 205.380 109.980 205.550 ;
        RECT 111.245 204.055 111.415 215.345 ;
        RECT 98.885 203.885 111.415 204.055 ;
        RECT 100.800 188.815 101.700 189.000 ;
        RECT 98.885 188.645 111.415 188.815 ;
        RECT 98.885 177.355 99.055 188.645 ;
        RECT 100.800 188.400 101.700 188.645 ;
        RECT 100.800 187.420 101.700 187.500 ;
        RECT 100.380 187.250 109.980 187.420 ;
        RECT 100.380 178.850 100.550 187.250 ;
        RECT 100.800 187.200 101.700 187.250 ;
        RECT 101.180 186.740 109.180 186.910 ;
        RECT 100.950 179.530 101.120 186.570 ;
        RECT 109.240 179.530 109.410 186.570 ;
        RECT 101.180 179.190 109.180 179.360 ;
        RECT 109.810 178.850 109.980 187.250 ;
        RECT 100.380 178.680 109.980 178.850 ;
        RECT 111.245 177.355 111.415 188.645 ;
        RECT 98.885 177.185 111.415 177.355 ;
        RECT 98.885 161.345 111.415 161.515 ;
        RECT 98.885 150.055 99.055 161.345 ;
        RECT 100.800 160.120 101.700 160.200 ;
        RECT 100.380 159.950 109.980 160.120 ;
        RECT 100.380 151.550 100.550 159.950 ;
        RECT 100.800 159.900 101.700 159.950 ;
        RECT 101.180 159.440 109.180 159.610 ;
        RECT 100.950 152.230 101.120 159.270 ;
        RECT 109.240 152.230 109.410 159.270 ;
        RECT 101.180 151.890 109.180 152.060 ;
        RECT 109.810 151.550 109.980 159.950 ;
        RECT 100.380 151.380 109.980 151.550 ;
        RECT 111.245 150.055 111.415 161.345 ;
        RECT 98.885 149.885 111.415 150.055 ;
        RECT 108.900 143.515 109.800 143.700 ;
        RECT 98.885 143.345 111.415 143.515 ;
        RECT 98.885 132.055 99.055 143.345 ;
        RECT 108.900 143.100 109.800 143.345 ;
        RECT 108.900 142.120 109.500 142.200 ;
        RECT 100.380 141.950 109.980 142.120 ;
        RECT 100.380 133.550 100.550 141.950 ;
        RECT 108.900 141.900 109.500 141.950 ;
        RECT 101.180 141.440 109.180 141.610 ;
        RECT 100.950 134.230 101.120 141.270 ;
        RECT 109.240 134.230 109.410 141.270 ;
        RECT 101.180 133.890 109.180 134.060 ;
        RECT 109.810 133.550 109.980 141.950 ;
        RECT 100.380 133.380 109.980 133.550 ;
        RECT 111.245 132.055 111.415 143.345 ;
        RECT 98.885 131.885 111.415 132.055 ;
        RECT 106.730 60.560 149.050 60.730 ;
        RECT 106.730 7.900 106.900 60.560 ;
        RECT 107.380 8.380 107.730 10.540 ;
        RECT 148.050 8.380 148.400 10.540 ;
        RECT 147.000 7.900 147.600 8.100 ;
        RECT 148.880 7.900 149.050 60.560 ;
        RECT 106.730 7.730 149.050 7.900 ;
        RECT 149.830 60.640 158.950 60.810 ;
        RECT 149.830 7.900 150.000 60.640 ;
        RECT 150.480 8.380 150.830 10.540 ;
        RECT 157.950 9.000 158.300 10.540 ;
        RECT 157.800 8.400 158.400 9.000 ;
        RECT 157.950 8.380 158.300 8.400 ;
        RECT 157.800 7.900 158.400 8.100 ;
        RECT 158.780 7.900 158.950 60.640 ;
        RECT 149.830 7.730 158.950 7.900 ;
        RECT 147.000 7.500 147.600 7.730 ;
        RECT 157.800 7.500 158.400 7.730 ;
      LAYER mcon ;
        RECT 152.560 222.340 152.850 222.510 ;
        RECT 151.680 221.400 151.850 221.700 ;
        RECT 152.250 221.210 152.420 222.090 ;
        RECT 152.990 221.210 153.160 222.090 ;
        RECT 152.560 220.790 152.850 220.960 ;
        RECT 155.060 222.330 155.350 222.500 ;
        RECT 154.750 220.655 154.920 222.035 ;
        RECT 155.490 220.655 155.660 222.035 ;
        RECT 156.060 221.510 156.230 221.780 ;
        RECT 155.060 220.190 155.350 220.360 ;
        RECT 152.560 218.650 152.850 218.820 ;
        RECT 151.680 218.100 151.850 218.400 ;
        RECT 152.250 217.520 152.420 218.400 ;
        RECT 152.990 217.520 153.160 218.400 ;
        RECT 152.560 217.100 152.850 217.270 ;
        RECT 155.060 218.640 155.350 218.810 ;
        RECT 154.750 216.965 154.920 218.345 ;
        RECT 155.490 216.965 155.660 218.345 ;
        RECT 156.060 217.710 156.230 217.980 ;
        RECT 155.060 216.500 155.350 216.670 ;
        RECT 100.200 215.400 101.400 215.700 ;
        RECT 101.260 213.440 109.100 213.610 ;
        RECT 100.950 206.310 101.120 213.190 ;
        RECT 109.240 206.310 109.410 213.190 ;
        RECT 101.260 205.890 109.100 206.060 ;
        RECT 101.260 186.740 109.100 186.910 ;
        RECT 100.950 179.610 101.120 186.490 ;
        RECT 109.240 179.610 109.410 186.490 ;
        RECT 101.260 179.190 109.100 179.360 ;
        RECT 101.260 159.440 109.100 159.610 ;
        RECT 100.950 152.310 101.120 159.190 ;
        RECT 109.240 152.310 109.410 159.190 ;
        RECT 101.260 151.890 109.100 152.060 ;
        RECT 101.260 141.440 109.100 141.610 ;
        RECT 100.950 134.310 101.120 141.190 ;
        RECT 109.240 134.310 109.410 141.190 ;
        RECT 101.260 133.890 109.100 134.060 ;
        RECT 107.400 8.400 107.700 10.200 ;
        RECT 157.800 8.400 158.400 9.000 ;
      LAYER met1 ;
        RECT 152.500 222.530 155.400 222.600 ;
        RECT 152.500 222.300 155.410 222.530 ;
        RECT 151.650 221.700 151.880 221.760 ;
        RECT 152.220 221.700 152.450 222.150 ;
        RECT 152.960 221.800 153.190 222.150 ;
        RECT 154.720 221.800 154.950 222.095 ;
        RECT 155.460 221.800 155.690 222.095 ;
        RECT 156.000 221.800 156.300 222.600 ;
        RECT 145.750 221.400 152.450 221.700 ;
        RECT 152.900 221.500 155.000 221.800 ;
        RECT 155.460 221.500 156.300 221.800 ;
        RECT 151.650 221.340 151.880 221.400 ;
        RECT 152.220 221.150 152.450 221.400 ;
        RECT 152.960 221.150 153.190 221.500 ;
        RECT 152.500 220.760 152.910 220.990 ;
        RECT 153.800 219.900 154.100 221.500 ;
        RECT 154.720 220.595 154.950 221.500 ;
        RECT 155.460 220.595 155.690 221.500 ;
        RECT 155.000 220.160 155.410 220.390 ;
        RECT 153.750 219.600 154.150 219.900 ;
        RECT 153.800 218.900 154.100 219.600 ;
        RECT 152.400 218.600 155.500 218.900 ;
        RECT 151.650 218.400 151.880 218.460 ;
        RECT 152.220 218.400 152.450 218.460 ;
        RECT 145.750 218.100 152.450 218.400 ;
        RECT 151.650 218.040 151.880 218.100 ;
        RECT 152.220 217.460 152.450 218.100 ;
        RECT 152.960 218.000 153.190 218.460 ;
        RECT 154.720 218.000 154.950 218.405 ;
        RECT 152.960 217.700 154.950 218.000 ;
        RECT 152.960 217.460 153.190 217.700 ;
        RECT 100.150 216.300 101.450 217.200 ;
        RECT 152.500 217.070 152.910 217.300 ;
        RECT 100.200 215.730 101.400 216.300 ;
        RECT 100.140 215.370 101.460 215.730 ;
        RECT 153.400 215.700 153.700 217.700 ;
        RECT 154.720 216.905 154.950 217.700 ;
        RECT 155.460 218.000 155.690 218.405 ;
        RECT 156.000 218.000 156.300 221.500 ;
        RECT 155.460 217.700 156.300 218.000 ;
        RECT 155.460 216.905 155.690 217.700 ;
        RECT 156.000 217.000 156.300 217.700 ;
        RECT 155.000 216.470 155.410 216.700 ;
        RECT 155.950 216.400 156.350 217.000 ;
        RECT 100.200 214.230 101.400 215.370 ;
        RECT 153.250 214.800 153.950 215.700 ;
        RECT 100.200 213.870 101.460 214.230 ;
        RECT 100.200 213.640 101.400 213.870 ;
        RECT 100.200 213.410 109.160 213.640 ;
        RECT 100.200 212.700 101.400 213.410 ;
        RECT 100.920 206.250 101.150 212.700 ;
        RECT 109.210 211.500 109.440 213.250 ;
        RECT 109.200 210.600 112.550 211.500 ;
        RECT 109.210 206.250 109.440 210.600 ;
        RECT 101.200 205.860 109.160 206.090 ;
        RECT 100.750 189.300 101.750 190.200 ;
        RECT 100.800 189.030 101.700 189.300 ;
        RECT 100.740 188.370 101.760 189.030 ;
        RECT 100.800 187.530 101.700 188.370 ;
        RECT 100.740 187.170 101.760 187.530 ;
        RECT 100.800 186.940 101.700 187.170 ;
        RECT 100.800 186.710 109.160 186.940 ;
        RECT 100.800 185.700 101.700 186.710 ;
        RECT 100.920 179.550 101.150 185.700 ;
        RECT 109.210 183.300 109.440 186.550 ;
        RECT 109.200 182.400 112.550 183.300 ;
        RECT 109.210 179.550 109.440 182.400 ;
        RECT 101.200 179.160 109.160 179.390 ;
        RECT 100.750 162.000 101.750 162.900 ;
        RECT 100.800 160.230 101.700 162.000 ;
        RECT 100.740 159.870 101.760 160.230 ;
        RECT 100.800 159.640 101.700 159.870 ;
        RECT 100.800 159.410 109.160 159.640 ;
        RECT 100.800 158.400 101.700 159.410 ;
        RECT 100.920 152.250 101.150 158.400 ;
        RECT 109.210 156.300 109.440 159.250 ;
        RECT 109.200 155.400 112.850 156.300 ;
        RECT 109.210 152.250 109.440 155.400 ;
        RECT 101.200 151.860 109.160 152.090 ;
        RECT 108.850 144.000 109.850 144.900 ;
        RECT 108.900 143.730 109.800 144.000 ;
        RECT 108.840 143.070 109.860 143.730 ;
        RECT 108.900 142.230 109.800 143.070 ;
        RECT 108.840 141.870 109.800 142.230 ;
        RECT 108.900 141.640 109.800 141.870 ;
        RECT 101.200 141.410 109.800 141.640 ;
        RECT 100.920 141.000 101.150 141.250 ;
        RECT 96.900 140.700 101.150 141.000 ;
        RECT 96.850 139.500 101.150 140.700 ;
        RECT 108.900 140.400 109.800 141.410 ;
        RECT 96.900 138.300 101.150 139.500 ;
        RECT 96.850 137.100 101.150 138.300 ;
        RECT 96.900 135.900 101.150 137.100 ;
        RECT 96.850 134.700 101.150 135.900 ;
        RECT 96.900 134.400 101.150 134.700 ;
        RECT 100.920 134.250 101.150 134.400 ;
        RECT 109.210 134.250 109.440 140.400 ;
        RECT 101.200 133.860 109.160 134.090 ;
        RECT 103.800 10.260 107.700 10.500 ;
        RECT 103.800 8.400 107.730 10.260 ;
        RECT 107.370 8.340 107.730 8.400 ;
        RECT 148.020 8.780 148.430 8.840 ;
        RECT 150.450 8.780 150.860 8.840 ;
        RECT 148.020 8.380 150.860 8.780 ;
        RECT 148.020 8.320 148.430 8.380 ;
        RECT 150.450 8.320 150.860 8.380 ;
        RECT 157.740 8.370 158.460 9.030 ;
        RECT 157.800 8.130 158.400 8.370 ;
        RECT 146.940 7.470 147.660 8.130 ;
        RECT 157.740 7.470 158.460 8.130 ;
        RECT 147.000 5.700 147.600 7.470 ;
        RECT 157.800 5.700 158.400 7.470 ;
        RECT 146.950 5.100 147.650 5.700 ;
        RECT 157.750 5.100 158.450 5.700 ;
      LAYER via ;
        RECT 153.800 222.300 154.100 222.600 ;
        RECT 145.800 221.400 146.700 221.700 ;
        RECT 153.800 219.600 154.100 219.900 ;
        RECT 145.800 218.100 146.700 218.400 ;
        RECT 100.200 216.300 101.400 217.200 ;
        RECT 156.000 216.400 156.300 217.000 ;
        RECT 153.300 214.800 153.900 215.700 ;
        RECT 111.600 210.600 112.500 211.500 ;
        RECT 100.800 189.300 101.700 190.200 ;
        RECT 111.600 182.400 112.500 183.300 ;
        RECT 100.800 162.000 101.700 162.900 ;
        RECT 111.900 155.400 112.800 156.300 ;
        RECT 108.900 144.000 109.800 144.900 ;
        RECT 96.900 139.500 98.100 140.700 ;
        RECT 96.900 137.100 98.100 138.300 ;
        RECT 96.900 134.700 98.100 135.900 ;
        RECT 104.100 8.700 106.200 10.200 ;
        RECT 148.860 8.390 149.460 8.760 ;
        RECT 147.000 5.100 147.600 5.700 ;
        RECT 157.800 5.100 158.400 5.700 ;
      LAYER met2 ;
        RECT 153.800 222.250 154.100 224.750 ;
        RECT 145.800 221.350 146.700 221.750 ;
        RECT 139.500 219.900 140.100 219.950 ;
        RECT 153.800 219.900 154.100 219.950 ;
        RECT 139.500 219.300 154.200 219.900 ;
        RECT 139.500 219.250 140.100 219.300 ;
        RECT 145.800 218.050 146.700 218.450 ;
        RECT 100.200 216.250 101.400 217.250 ;
        RECT 100.800 190.200 101.700 190.250 ;
        RECT 111.600 190.200 112.500 211.550 ;
        RECT 100.800 189.300 112.500 190.200 ;
        RECT 100.800 189.250 101.700 189.300 ;
        RECT 111.600 189.000 112.500 189.300 ;
        RECT 100.800 162.900 101.700 162.950 ;
        RECT 111.600 162.900 112.500 183.350 ;
        RECT 100.800 162.000 112.500 162.900 ;
        RECT 100.800 161.950 101.700 162.000 ;
        RECT 147.900 159.550 148.500 219.300 ;
        RECT 156.000 216.350 156.300 217.050 ;
        RECT 153.300 214.750 153.900 215.750 ;
        RECT 108.900 144.900 109.800 144.950 ;
        RECT 111.900 144.900 112.800 156.350 ;
        RECT 108.900 144.000 112.800 144.900 ;
        RECT 108.900 143.950 109.800 144.000 ;
        RECT 96.900 139.450 98.100 140.750 ;
        RECT 96.900 137.050 98.100 138.350 ;
        RECT 96.900 134.650 98.100 135.950 ;
        RECT 104.100 8.650 106.200 10.250 ;
        RECT 148.860 8.340 149.460 8.810 ;
        RECT 49.500 5.700 50.100 5.750 ;
        RECT 147.000 5.700 147.600 5.750 ;
        RECT 157.800 5.700 158.400 5.750 ;
        RECT 49.500 5.100 158.400 5.700 ;
        RECT 49.500 5.050 50.100 5.100 ;
        RECT 147.000 5.050 147.600 5.100 ;
        RECT 157.800 5.050 158.400 5.100 ;
      LAYER via2 ;
        RECT 153.800 224.300 154.100 224.700 ;
        RECT 145.800 221.400 146.700 221.700 ;
        RECT 145.800 218.100 146.700 218.400 ;
        RECT 100.200 216.300 101.400 217.200 ;
        RECT 111.600 210.600 112.500 211.500 ;
        RECT 111.600 182.400 112.500 183.300 ;
        RECT 156.000 216.400 156.300 217.000 ;
        RECT 153.300 214.800 153.900 215.700 ;
        RECT 147.900 159.600 148.500 160.200 ;
        RECT 111.900 155.400 112.800 156.300 ;
        RECT 96.900 139.500 98.100 140.700 ;
        RECT 96.900 137.100 98.100 138.300 ;
        RECT 96.900 134.700 98.100 135.900 ;
        RECT 104.100 8.700 106.200 10.200 ;
        RECT 148.860 8.390 149.460 8.760 ;
      LAYER met3 ;
        RECT 153.750 224.700 154.150 224.725 ;
        RECT 153.650 224.300 154.250 224.700 ;
        RECT 153.750 224.275 154.150 224.300 ;
        RECT 145.450 222.500 147.050 224.000 ;
        RECT 139.450 219.275 140.150 219.925 ;
        RECT 145.500 218.000 147.000 222.500 ;
        RECT 100.150 217.200 101.450 217.225 ;
        RECT 100.150 217.000 143.750 217.200 ;
        RECT 155.950 217.000 156.350 217.025 ;
        RECT 100.150 216.400 156.350 217.000 ;
        RECT 100.150 216.300 143.750 216.400 ;
        RECT 155.950 216.375 156.350 216.400 ;
        RECT 100.150 216.275 101.450 216.300 ;
        RECT 111.550 210.575 112.550 211.525 ;
        RECT 113.500 189.500 139.995 215.500 ;
        RECT 153.250 214.775 153.950 215.725 ;
        RECT 111.550 182.375 112.550 183.325 ;
        RECT 113.400 162.300 139.895 188.300 ;
        RECT 153.300 187.200 153.900 214.775 ;
        RECT 140.350 186.600 153.900 187.200 ;
        RECT 111.850 155.375 112.850 156.325 ;
        RECT 64.200 119.700 95.695 145.700 ;
        RECT 96.900 140.725 98.100 141.000 ;
        RECT 96.850 139.475 98.150 140.725 ;
        RECT 96.900 138.325 98.100 139.475 ;
        RECT 96.850 137.075 98.150 138.325 ;
        RECT 96.900 135.925 98.100 137.075 ;
        RECT 96.850 134.675 98.150 135.925 ;
        RECT 113.400 135.000 139.895 161.000 ;
        RECT 147.850 160.200 148.550 160.225 ;
        RECT 140.350 159.600 148.550 160.200 ;
        RECT 147.850 159.575 148.550 159.600 ;
        RECT 96.900 10.500 98.100 134.675 ;
        RECT 96.900 8.400 106.500 10.500 ;
        RECT 148.810 8.365 149.510 8.785 ;
        RECT 49.450 5.075 50.150 5.725 ;
      LAYER via3 ;
        RECT 153.700 224.300 154.200 224.700 ;
        RECT 145.500 222.500 147.000 224.000 ;
        RECT 139.500 219.300 140.100 219.900 ;
        RECT 142.200 216.300 143.700 217.200 ;
        RECT 111.600 210.600 112.500 211.500 ;
        RECT 139.575 189.640 139.895 215.360 ;
        RECT 111.600 182.400 112.500 183.300 ;
        RECT 139.475 162.440 139.795 188.160 ;
        RECT 140.400 186.600 141.300 187.200 ;
        RECT 111.900 155.400 112.800 156.300 ;
        RECT 95.275 119.840 95.595 145.560 ;
        RECT 96.900 139.500 98.100 140.700 ;
        RECT 96.900 137.100 98.100 138.300 ;
        RECT 96.900 134.700 98.100 135.900 ;
        RECT 139.475 135.140 139.795 160.860 ;
        RECT 140.400 159.600 141.300 160.200 ;
        RECT 148.860 8.390 149.460 8.760 ;
        RECT 49.500 5.100 50.100 5.700 ;
      LAYER met4 ;
        RECT 4.290 224.760 4.295 225.760 ;
        RECT 3.995 224.005 4.295 224.760 ;
        RECT 7.670 224.005 7.970 224.760 ;
        RECT 11.350 224.005 11.650 224.760 ;
        RECT 15.030 224.005 15.330 224.760 ;
        RECT 18.710 224.005 19.010 224.760 ;
        RECT 22.390 224.005 22.690 224.760 ;
        RECT 26.070 224.005 26.370 224.760 ;
        RECT 29.750 224.005 30.050 224.760 ;
        RECT 33.430 224.005 33.730 224.760 ;
        RECT 37.110 224.005 37.410 224.760 ;
        RECT 40.790 224.005 41.090 224.760 ;
        RECT 44.470 224.005 44.770 224.760 ;
        RECT 48.150 224.005 48.450 224.760 ;
        RECT 51.830 224.005 52.130 224.760 ;
        RECT 55.510 224.005 55.810 224.760 ;
        RECT 59.190 224.005 59.490 224.760 ;
        RECT 62.870 224.005 63.170 224.760 ;
        RECT 66.550 224.005 66.850 224.760 ;
        RECT 70.230 224.005 70.530 224.760 ;
        RECT 73.910 224.005 74.210 224.760 ;
        RECT 77.590 224.005 77.890 224.760 ;
        RECT 81.270 224.005 81.570 224.760 ;
        RECT 84.950 224.005 85.250 224.760 ;
        RECT 88.630 224.005 88.930 224.760 ;
        RECT 153.695 224.650 154.205 224.705 ;
        RECT 154.870 224.650 155.170 224.760 ;
        RECT 153.695 224.350 155.170 224.650 ;
        RECT 153.695 224.295 154.205 224.350 ;
        RECT 3.995 224.000 88.945 224.005 ;
        RECT 145.495 224.000 147.005 224.005 ;
        RECT 3.995 223.705 147.005 224.000 ;
        RECT 4.000 223.500 147.005 223.705 ;
        RECT 49.000 222.500 147.005 223.500 ;
        RECT 49.000 220.760 50.500 222.500 ;
        RECT 145.495 222.495 147.005 222.500 ;
        RECT 139.495 219.295 140.105 219.905 ;
        RECT 139.500 215.440 140.100 219.295 ;
        RECT 142.195 216.295 142.200 217.205 ;
        RECT 143.700 216.295 143.705 217.205 ;
        RECT 139.495 215.100 140.100 215.440 ;
        RECT 111.595 211.500 112.505 211.505 ;
        RECT 114.195 211.500 138.805 214.805 ;
        RECT 111.595 210.600 138.805 211.500 ;
        RECT 111.595 210.595 112.505 210.600 ;
        RECT 114.195 190.195 138.805 210.600 ;
        RECT 139.495 189.560 139.975 215.100 ;
        RECT 139.395 188.100 139.875 188.240 ;
        RECT 111.595 183.300 112.505 183.305 ;
        RECT 114.095 183.300 138.705 187.605 ;
        RECT 111.595 182.400 138.705 183.300 ;
        RECT 111.595 182.395 112.505 182.400 ;
        RECT 114.095 162.995 138.705 182.400 ;
        RECT 139.395 186.000 141.600 188.100 ;
        RECT 139.395 162.360 139.875 186.000 ;
        RECT 139.395 160.800 139.875 160.940 ;
        RECT 111.895 156.300 112.805 156.305 ;
        RECT 114.095 156.300 138.705 160.305 ;
        RECT 111.895 155.400 138.705 156.300 ;
        RECT 111.895 155.395 112.805 155.400 ;
        RECT 64.895 139.200 94.505 145.005 ;
        RECT 95.195 141.000 95.675 145.640 ;
        RECT 50.500 128.400 94.505 139.200 ;
        RECT 95.100 140.705 98.100 141.000 ;
        RECT 95.100 139.495 98.105 140.705 ;
        RECT 95.100 138.305 98.100 139.495 ;
        RECT 95.100 137.095 98.105 138.305 ;
        RECT 95.100 135.905 98.100 137.095 ;
        RECT 95.100 134.695 98.105 135.905 ;
        RECT 114.095 135.695 138.705 155.400 ;
        RECT 139.395 159.000 141.600 160.800 ;
        RECT 139.395 135.060 139.875 159.000 ;
        RECT 95.100 134.400 98.100 134.695 ;
        RECT 64.895 120.395 94.505 128.400 ;
        RECT 95.195 119.760 95.675 134.400 ;
        RECT 148.850 8.765 149.450 8.790 ;
        RECT 148.850 8.385 149.465 8.765 ;
        RECT 148.850 7.250 149.450 8.385 ;
        RECT 148.850 6.650 157.160 7.250 ;
        RECT 156.560 1.000 157.160 6.650 ;
  END
END tt_um_urish_charge_pump
END LIBRARY

