magic
tech sky130A
magscale 1 2
timestamp 1711870259
<< metal3 >>
rect -3150 2572 3149 2600
rect -3150 -2572 3065 2572
rect 3129 -2572 3149 2572
rect -3150 -2600 3149 -2572
<< via3 >>
rect 3065 -2572 3129 2572
<< mimcap >>
rect -3050 2460 2950 2500
rect -3050 -2460 -3010 2460
rect 2910 -2460 2950 2460
rect -3050 -2500 2950 -2460
<< mimcapcontact >>
rect -3010 -2460 2910 2460
<< metal4 >>
rect 3049 2572 3145 2588
rect -3011 2460 2911 2461
rect -3011 -2460 -3010 2460
rect 2910 -2460 2911 2460
rect -3011 -2461 2911 -2460
rect 3049 -2572 3065 2572
rect 3129 -2572 3145 2572
rect 3049 -2588 3145 -2572
<< properties >>
string FIXED_BBOX -3150 -2600 3050 2600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 25.0 val 1.52k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
