* NGSPICE file created from tt_um_urish_charge_pump.ext - technology: sky130A

.subckt tt_um_urish_charge_pump clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VPWR VGND
X0 clka clk.t0 VGND.t5 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.45
X1 stage2.t4 clkb.t2 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X2 stage3.t3 stage2.t1 stage2.t3 stage2.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X3 VGND.t4 ua[0].t1 VGND.t3 sky130_fd_pr__res_xhigh_po_0p35 l=493.37
X4 VGND.t6 vout sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X5 stage3.t4 clka.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X6 clkb.t1 clka VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.45
X7 VPWR.t5 clk.t1 clka VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.45
X8 stage3.t2 stage3.t0 vout stage3.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X9 stage2.t0 stage1.t1 stage1.t3 stage1.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X10 ua[0].t0 vout VGND.t2 sky130_fd_pr__res_xhigh_po_0p35 l=2.45857k
X11 stage1.t0 VPWR.t2 VPWR.t4 VPWR.t3 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X12 stage1.t4 clka.t1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X13 VPWR.t1 clka.t2 clkb.t0 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.45
R0 clk.n0 clk.t1 276.433
R1 clk.n0 clk.t0 244.831
R2 clk clk.n0 12.3379
R3 VGND.n70 VGND.n4 54934
R4 VGND.n70 VGND.n5 54934
R5 VGND.n71 VGND.n4 54934
R6 VGND.n71 VGND.n5 54934
R7 VGND.n15 VGND.n6 35743.9
R8 VGND.n10 VGND.n7 35743.9
R9 VGND.n15 VGND.n7 35743.9
R10 VGND.n67 VGND.n18 18300
R11 VGND.n67 VGND.n66 8364.42
R12 VGND.n68 VGND.n67 4592.88
R13 VGND.n72 VGND.n3 3569.32
R14 VGND.n69 VGND.n3 3569.32
R15 VGND.n69 VGND.n2 3569.32
R16 VGND.n23 VGND.n20 2479.88
R17 VGND.n65 VGND.n20 2479.88
R18 VGND.n23 VGND.n21 2479.88
R19 VGND.n65 VGND.n21 2479.88
R20 VGND.n54 VGND.n19 2479.88
R21 VGND.n56 VGND.n19 2479.88
R22 VGND.n56 VGND.n55 2479.88
R23 VGND.n55 VGND.n54 2479.88
R24 VGND.n11 VGND.n8 2322.45
R25 VGND.n14 VGND.n8 2322.45
R26 VGND.n14 VGND.n13 2322.45
R27 VGND.n73 VGND.n2 2091.67
R28 VGND.n12 VGND.n11 2026.92
R29 VGND.n73 VGND.n72 1445.27
R30 VGND.t0 VGND.n18 415.678
R31 VGND.n66 VGND.t0 415.678
R32 VGND.n13 VGND.n12 263.154
R33 VGND.n25 VGND.n21 195
R34 VGND.n21 VGND.t0 195
R35 VGND.n22 VGND.n20 195
R36 VGND.n20 VGND.t0 195
R37 VGND.n54 VGND.n52 195
R38 VGND.n54 VGND.t0 195
R39 VGND.n57 VGND.n56 195
R40 VGND.n56 VGND.t0 195
R41 VGND.n24 VGND.n22 161.13
R42 VGND.n64 VGND.n22 161.13
R43 VGND.n25 VGND.n24 161.13
R44 VGND.n53 VGND.n52 161.13
R45 VGND.n57 VGND.n53 161.13
R46 VGND.n58 VGND.n57 161.13
R47 VGND.n63 VGND.n25 153.601
R48 VGND.n59 VGND.n52 139.294
R49 VGND.n65 VGND.n64 117.001
R50 VGND.n66 VGND.n65 117.001
R51 VGND.n24 VGND.n23 117.001
R52 VGND.n23 VGND.n18 117.001
R53 VGND.n55 VGND.n53 117.001
R54 VGND.n55 VGND.n18 117.001
R55 VGND.n58 VGND.n19 117.001
R56 VGND.n66 VGND.n19 117.001
R57 VGND.n60 VGND.t1 84.0308
R58 VGND.n62 VGND.t5 83.9547
R59 VGND.n17 VGND.n16 31.7634
R60 VGND.n10 VGND.n9 28.5239
R61 VGND.n75 VGND.n74 27.133
R62 VGND.n16 VGND.t3 24.7421
R63 VGND.t2 VGND.n17 24.7421
R64 VGND.n13 VGND.n7 24.3755
R65 VGND.n7 VGND.t3 24.3755
R66 VGND.n8 VGND.n6 24.3755
R67 VGND.n9 VGND.n6 24.34
R68 VGND.n59 VGND.n58 21.8358
R69 VGND.n68 VGND.n5 18.8551
R70 VGND.t2 VGND.n68 9.64362
R71 VGND.n63 VGND.n62 9.3005
R72 VGND.n60 VGND.n59 9.3005
R73 VGND.n64 VGND.n63 7.52991
R74 VGND.n61 VGND.n60 5.60682
R75 VGND.n62 VGND.n61 5.50342
R76 VGND.n1 VGND.t4 4.88866
R77 VGND.n72 VGND.n71 4.79558
R78 VGND.n71 VGND.t2 4.79558
R79 VGND.n70 VGND.n69 4.79558
R80 VGND.t2 VGND.n70 4.79558
R81 VGND.n39 VGND 4.20543
R82 VGND.n74 VGND.n73 3.93011
R83 VGND.n74 VGND.n1 3.85511
R84 VGND.n76 VGND.n75 3.8545
R85 VGND.n15 VGND.n14 3.82403
R86 VGND.n16 VGND.n15 3.82403
R87 VGND.n11 VGND.n10 3.82403
R88 VGND.n5 VGND.n3 3.82403
R89 VGND.n4 VGND.n2 3.82403
R90 VGND.n17 VGND.n4 3.82403
R91 VGND.n40 VGND.n39 2.61057
R92 VGND.n12 VGND.n1 2.3255
R93 VGND.n61 VGND.n51 2.23174
R94 VGND.n26 uio_oe[7] 1.43262
R95 VGND.n27 VGND.n26 0.438736
R96 VGND VGND.n76 0.365382
R97 VGND.n38 VGND.n37 0.342995
R98 VGND.n37 VGND.n36 0.342995
R99 VGND.n36 VGND.n35 0.342995
R100 VGND.n35 VGND.n34 0.342995
R101 VGND.n34 VGND.n33 0.342995
R102 VGND.n33 VGND.n32 0.342995
R103 VGND.n32 VGND.n31 0.342995
R104 VGND.n31 VGND.n30 0.342995
R105 VGND.n30 VGND.n29 0.342995
R106 VGND.n29 VGND.n28 0.342995
R107 VGND.n28 VGND.n27 0.342995
R108 VGND.n38 uio_out[3] 0.118783
R109 VGND.n37 uio_out[4] 0.118783
R110 VGND.n36 uio_out[5] 0.118783
R111 VGND.n35 uio_out[6] 0.118783
R112 VGND.n34 uio_out[7] 0.118783
R113 VGND.n33 uio_oe[0] 0.118783
R114 VGND.n32 uio_oe[1] 0.118783
R115 VGND.n31 uio_oe[2] 0.118783
R116 VGND.n30 uio_oe[3] 0.118783
R117 VGND.n29 uio_oe[4] 0.118783
R118 VGND.n28 uio_oe[5] 0.118783
R119 VGND.n27 uio_oe[6] 0.118783
R120 VGND.n51 uo_out[0] 0.118783
R121 VGND.n50 uo_out[1] 0.118783
R122 VGND.n49 uo_out[2] 0.118783
R123 VGND.n48 uo_out[3] 0.118783
R124 VGND.n47 uo_out[4] 0.118783
R125 VGND.n46 uo_out[5] 0.118783
R126 VGND.n45 uo_out[6] 0.118783
R127 VGND.n44 uo_out[7] 0.118783
R128 VGND.n43 uio_out[0] 0.118783
R129 VGND.n42 uio_out[1] 0.118783
R130 VGND.n41 uio_out[2] 0.118783
R131 VGND.n51 VGND.n50 0.115424
R132 VGND.n50 VGND.n49 0.115424
R133 VGND.n49 VGND.n48 0.115424
R134 VGND.n48 VGND.n47 0.115424
R135 VGND.n47 VGND.n46 0.115424
R136 VGND.n46 VGND.n45 0.115424
R137 VGND.n45 VGND.n44 0.115424
R138 VGND.n44 VGND.n43 0.115424
R139 VGND.n43 VGND.n42 0.115424
R140 VGND.n42 VGND.n41 0.115424
R141 VGND.n40 VGND.n38 0.0890704
R142 VGND.n41 VGND.n40 0.0701412
R143 VGND.n0 VGND.t6 0.0297714
R144 VGND.n26 uio_oe[7] 0.0252647
R145 VGND.n9 VGND.t3 0.0204508
R146 VGND.n39 VGND.n0 0.0164673
R147 VGND.n76 VGND.n0 0.0164673
R148 VGND.n75 VGND 0.0130333
R149 clka clka.t2 276.433
R150 clka.n0 clka.t0 19.2376
R151 clka.n0 clka.t1 10.2333
R152 clka clka.n0 6.03696
R153 stage2.n7 stage2.n2 10330.9
R154 stage2.n6 stage2.n5 10330.9
R155 stage2.n5 stage2.t2 1841.91
R156 stage2.n7 stage2.n3 1841.91
R157 stage2.n8 stage2.n1 671.247
R158 stage2.n4 stage2.n1 671.247
R159 stage2.n4 stage2.n0 671.247
R160 stage2.t3 stage2.n8 360.659
R161 stage2.t3 stage2.n0 281.224
R162 stage2.t3 stage2.t1 31.6676
R163 stage2.n8 stage2.n7 25.4353
R164 stage2.n5 stage2.n4 25.4353
R165 stage2.n6 stage2.n1 23.4005
R166 stage2.n2 stage2.n0 23.4005
R167 stage2.t2 stage2.n2 19.1855
R168 stage2.n3 stage2.n6 19.1855
R169 stage2.t4 stage2.t0 13.1042
R170 stage2.n3 stage2.t2 8.34551
R171 stage2.t3 stage2.t4 8.27133
R172 clkb clkb.t0 167.643
R173 clkb clkb.t1 83.7335
R174 clkb clkb.t2 9.32862
R175 stage3.n8 stage3.n3 10330.9
R176 stage3.n7 stage3.n4 10330.9
R177 stage3.n19 stage3.n18 6978.85
R178 stage3.n18 stage3.n17 6978.85
R179 stage3.n17 stage3.n14 6978.85
R180 stage3.n19 stage3.n14 6978.85
R181 stage3.n20 stage3.n13 3802.7
R182 stage3.n16 stage3.n13 3802.7
R183 stage3.n16 stage3.n12 3802.7
R184 stage3.n20 stage3.n12 3802.7
R185 stage3.t1 stage3.n3 1841.91
R186 stage3.n5 stage3.n4 1841.91
R187 stage3.n21 stage3.n11 890.354
R188 stage3.n15 stage3.n11 890.354
R189 stage3.n15 stage3.n10 890.354
R190 stage3.n9 stage3.n2 671.247
R191 stage3.n6 stage3.n2 671.247
R192 stage3.n6 stage3.n1 671.247
R193 stage3.t4 stage3.n10 549.836
R194 stage3.n0 stage3.n1 358.776
R195 stage3.n0 stage3.n9 292.894
R196 stage3.t4 stage3.n21 291.954
R197 stage3.t4 stage3.t0 31.798
R198 stage3.n3 stage3.n2 25.4353
R199 stage3.n4 stage3.n1 25.4353
R200 stage3.n9 stage3.n8 23.4005
R201 stage3.n7 stage3.n6 23.4005
R202 stage3.n8 stage3.n5 19.1855
R203 stage3.t1 stage3.n7 19.1855
R204 stage3.t4 stage3.t2 13.8222
R205 stage3.t4 stage3.t3 13.743
R206 stage3.t4 stage3.n0 9.00675
R207 stage3.n5 stage3.t1 8.34551
R208 stage3.n13 stage3.n11 5.78175
R209 stage3.n18 stage3.n13 5.78175
R210 stage3.n12 stage3.n10 5.78175
R211 stage3.n14 stage3.n12 5.78175
R212 stage3.n21 stage3.n20 5.28621
R213 stage3.n20 stage3.n19 5.28621
R214 stage3.n16 stage3.n15 5.28621
R215 stage3.n17 stage3.n16 5.28621
R216 ua[0].n0 ua[0].t1 18.1143
R217 ua[0].n0 ua[0].t0 17.9393
R218 ua[0] ua[0].n0 10.2992
R219 VPWR.n32 VPWR.n26 10330.9
R220 VPWR.n30 VPWR.n29 10330.9
R221 VPWR.n43 VPWR.n40 6978.85
R222 VPWR.n45 VPWR.n40 6978.85
R223 VPWR.n44 VPWR.n43 6978.85
R224 VPWR.n45 VPWR.n44 6978.85
R225 VPWR.n42 VPWR.n38 3802.7
R226 VPWR.n46 VPWR.n38 3802.7
R227 VPWR.n42 VPWR.n39 3802.7
R228 VPWR.n46 VPWR.n39 3802.7
R229 VPWR.n29 VPWR.n28 1841.91
R230 VPWR.n32 VPWR.n31 1841.91
R231 VPWR.n16 VPWR.n5 1718.82
R232 VPWR.n12 VPWR.n5 1718.82
R233 VPWR.n16 VPWR.n6 1718.82
R234 VPWR.n12 VPWR.n6 1718.82
R235 VPWR.n10 VPWR.n3 1718.82
R236 VPWR.n10 VPWR.n4 1718.82
R237 VPWR.n18 VPWR.n4 1718.82
R238 VPWR.n18 VPWR.n3 1718.82
R239 VPWR.n47 VPWR.n37 890.354
R240 VPWR.n41 VPWR.n37 890.354
R241 VPWR.n41 VPWR.n36 890.354
R242 VPWR.n33 VPWR.n25 671.247
R243 VPWR.n27 VPWR.n25 671.247
R244 VPWR.n27 VPWR.n24 671.247
R245 VPWR.n48 VPWR.n47 539.282
R246 VPWR.n34 VPWR.n33 354.26
R247 VPWR.n48 VPWR.n36 303.988
R248 VPWR.n34 VPWR.n24 297.413
R249 VPWR.n13 VPWR.n8 183.341
R250 VPWR.n15 VPWR.n14 183.341
R251 VPWR.n14 VPWR.n13 183.341
R252 VPWR.n9 VPWR.n1 183.341
R253 VPWR.n9 VPWR.n2 183.341
R254 VPWR.n19 VPWR.n2 183.341
R255 VPWR.n20 VPWR.n1 169.036
R256 VPWR.n0 VPWR.t5 167.94
R257 VPWR.n21 VPWR.t1 167.881
R258 VPWR.n8 VPWR.n7 160.754
R259 VPWR.n17 VPWR.t0 121.004
R260 VPWR.n11 VPWR.t0 121.004
R261 VPWR.n14 VPWR.n6 61.6672
R262 VPWR.n6 VPWR.t0 61.6672
R263 VPWR.n8 VPWR.n5 61.6672
R264 VPWR.n5 VPWR.t0 61.6672
R265 VPWR.n3 VPWR.n1 61.6672
R266 VPWR.t0 VPWR.n3 61.6672
R267 VPWR.n4 VPWR.n2 61.6672
R268 VPWR.t0 VPWR.n4 61.6672
R269 VPWR.n23 VPWR.t2 31.8306
R270 VPWR.n13 VPWR.n12 26.4291
R271 VPWR.n12 VPWR.n11 26.4291
R272 VPWR.n16 VPWR.n15 26.4291
R273 VPWR.n17 VPWR.n16 26.4291
R274 VPWR.n10 VPWR.n9 26.4291
R275 VPWR.n11 VPWR.n10 26.4291
R276 VPWR.n19 VPWR.n18 26.4291
R277 VPWR.n18 VPWR.n17 26.4291
R278 VPWR.n33 VPWR.n32 25.4353
R279 VPWR.n29 VPWR.n27 25.4353
R280 VPWR.n30 VPWR.n25 23.4005
R281 VPWR.n26 VPWR.n24 23.4005
R282 VPWR.n15 VPWR.n7 22.5887
R283 VPWR.n28 VPWR.n26 19.1855
R284 VPWR.n31 VPWR.n30 19.1855
R285 VPWR.n20 VPWR.n19 14.3064
R286 VPWR.n23 VPWR.t4 13.9149
R287 VPWR.n7 VPWR.n0 9.3005
R288 VPWR.n21 VPWR.n20 9.3005
R289 VPWR VPWR.n50 7.20367
R290 VPWR.n50 VPWR.n22 7.05903
R291 VPWR.n47 VPWR.n46 5.78175
R292 VPWR.n46 VPWR.n45 5.78175
R293 VPWR.n42 VPWR.n41 5.78175
R294 VPWR.n43 VPWR.n42 5.78175
R295 VPWR.n39 VPWR.n37 5.28621
R296 VPWR.n44 VPWR.n39 5.28621
R297 VPWR.n38 VPWR.n36 5.28621
R298 VPWR.n40 VPWR.n38 5.28621
R299 VPWR.n35 VPWR.n34 4.6505
R300 VPWR.n31 VPWR.t3 4.17301
R301 VPWR.n28 VPWR.t3 4.17301
R302 VPWR.n50 VPWR.n49 3.42531
R303 VPWR.n49 VPWR.n48 3.1005
R304 VPWR.n22 VPWR.n0 1.46092
R305 VPWR.n49 VPWR.n35 0.15675
R306 VPWR.n35 VPWR.n23 0.0551875
R307 VPWR.n22 VPWR.n21 0.00258333
R308 stage1.n10 stage1.n4 10330.9
R309 stage1.n8 stage1.n7 10330.9
R310 stage1.n19 stage1.n16 6978.85
R311 stage1.n21 stage1.n16 6978.85
R312 stage1.n20 stage1.n19 6978.85
R313 stage1.n21 stage1.n20 6978.85
R314 stage1.n18 stage1.n14 3802.7
R315 stage1.n22 stage1.n14 3802.7
R316 stage1.n18 stage1.n15 3802.7
R317 stage1.n22 stage1.n15 3802.7
R318 stage1.n7 stage1.n6 1841.91
R319 stage1.n10 stage1.n9 1841.91
R320 stage1.n23 stage1.n13 890.354
R321 stage1.n17 stage1.n13 890.354
R322 stage1.n17 stage1.n12 890.354
R323 stage1.n11 stage1.n3 671.247
R324 stage1.n5 stage1.n3 671.247
R325 stage1.n5 stage1.n2 671.247
R326 stage1.n1 stage1.n23 572.424
R327 stage1.n0 stage1.n11 360.659
R328 stage1.n0 stage1.n2 281.224
R329 stage1.n1 stage1.n12 269.365
R330 stage1.n1 stage1.t1 31.6676
R331 stage1.n11 stage1.n10 25.4353
R332 stage1.n7 stage1.n5 25.4353
R333 stage1.n8 stage1.n3 23.4005
R334 stage1.n4 stage1.n2 23.4005
R335 stage1.n6 stage1.n4 19.1855
R336 stage1.n9 stage1.n8 19.1855
R337 stage1.n1 stage1.t3 13.8222
R338 stage1.t4 stage1.t0 13.5661
R339 stage1.n23 stage1.n22 5.78175
R340 stage1.n22 stage1.n21 5.78175
R341 stage1.n18 stage1.n17 5.78175
R342 stage1.n19 stage1.n18 5.78175
R343 stage1.n15 stage1.n13 5.28621
R344 stage1.n20 stage1.n15 5.28621
R345 stage1.n14 stage1.n12 5.28621
R346 stage1.n16 stage1.n14 5.28621
R347 stage1.n1 stage1.t4 5.03592
R348 stage1.n1 stage1.n0 4.91092
R349 stage1.n9 stage1.t2 4.17301
R350 stage1.n6 stage1.t2 4.17301
C0 ui_in[2] ui_in[1] 0.023797f
C1 VPWR uio_in[3] 1.03e-19
C2 rst_n clka 7.04e-19
C3 m2_3592_15598# m2_2584_17838# 0.151985f
C4 clka clkb 2.835f
C5 m2_2584_29654# m2_3592_27358# 0.091013f
C6 ui_in[5] ui_in[4] 0.023797f
C7 m2_2864_8934# m2_3648_12070# 0.135204f
C8 VPWR ui_in[1] 1.86e-20
C9 clk VPWR 0.418476f
C10 uio_in[0] uio_in[1] 0.023797f
C11 ui_in[0] VPWR 4.94e-20
C12 ui_in[6] VPWR 1.03e-19
C13 uio_in[0] ui_in[7] 0.023797f
C14 m2_1800_4342# m2_2864_8934# 0.00172f
C15 ui_in[3] ui_in[4] 0.023797f
C16 rst_n VPWR 4.94e-20
C17 VPWR clkb 1.72951f
C18 ua[0] VPWR 0.040036f
C19 uio_in[2] uio_in[3] 0.023797f
C20 ui_in[0] ui_in[1] 0.023797f
C21 VPWR uio_in[2] 1.03e-19
C22 VPWR uio_in[1] 1.03e-19
C23 ui_in[7] VPWR 1.03e-19
C24 VPWR ui_in[4] 1.03e-19
C25 rst_n clk 0.023797f
C26 uio_in[4] uio_in[3] 0.023797f
C27 clk clkb 0.001409f
C28 rst_n ui_in[0] 0.023797f
C29 uio_in[4] VPWR 1.03e-19
C30 ui_in[2] clka 3.03e-19
C31 uio_in[6] uio_in[5] 0.023797f
C32 uio_in[6] uio_in[7] 0.023797f
C33 m2_2864_23326# m2_3592_27358# 0.138713f
C34 ui_in[6] ui_in[7] 0.023797f
C35 ui_in[2] ui_in[3] 0.023797f
C36 m2_1800_4342# m2_3592_4230# 0.559432f
C37 ui_in[5] VPWR 1.03e-19
C38 m2_3592_42086# m2_3592_39062# 0.130452f
C39 m2_2472_13022# m2_3648_12070# 0.105624f
C40 clka VPWR 5.07751f
C41 m2_3592_35982# m2_2808_33406# 0.0711f
C42 m2_3592_35982# m2_3592_39062# 0.162853f
C43 m2_2472_13022# m2_2864_8934# 0.017782f
C44 uio_in[2] uio_in[1] 0.023797f
C45 clk ena 0.023797f
C46 ui_in[2] VPWR 1.03e-19
C47 uio_in[0] VPWR 1.03e-19
C48 dw_19800_30000# clka 0.101107f
C49 VPWR ui_in[3] 1.03e-19
C50 ui_in[6] ui_in[5] 0.023797f
C51 clka ui_in[1] 3.03e-19
C52 clk clka 0.275002f
C53 m2_2584_29654# m2_2808_33406# 0.041637f
C54 ui_in[0] clka 7.04e-19
C55 uio_in[4] uio_in[5] 0.023797f
C56 m2_3592_15598# m2_3648_12070# 0.104769f
C57 ua[1] VGND 0.123319f
C58 ua[2] VGND 0.123319f
C59 ua[3] VGND 0.123321f
C60 ua[4] VGND 0.123321f
C61 ua[5] VGND 0.122428f
C62 ua[6] VGND 0.122428f
C63 ua[7] VGND 0.122428f
C64 ena VGND 0.073297f
C65 rst_n VGND 0.048732f
C66 ui_in[0] VGND 0.048732f
C67 ui_in[1] VGND 0.05979f
C68 ui_in[2] VGND 0.05979f
C69 ui_in[3] VGND 0.05979f
C70 ui_in[4] VGND 0.05979f
C71 ui_in[5] VGND 0.05979f
C72 ui_in[6] VGND 0.05979f
C73 ui_in[7] VGND 0.05979f
C74 uio_in[0] VGND 0.05979f
C75 uio_in[1] VGND 0.05979f
C76 uio_in[2] VGND 0.05979f
C77 uio_in[3] VGND 0.05979f
C78 uio_in[4] VGND 0.05979f
C79 uio_in[5] VGND 0.05979f
C80 uio_in[6] VGND 0.05979f
C81 uio_in[7] VGND 0.083588f
C82 ua[0] VGND 2.69629f
C83 clk VGND 1.05257f
C84 VPWR VGND 49.875385f
C85 m2_3592_4230# VGND 2.41736f $ **FLOATING
C86 m2_1800_4342# VGND 11.662f $ **FLOATING
C87 m2_2864_8934# VGND 5.1283f $ **FLOATING
C88 m2_3648_12070# VGND 3.18023f $ **FLOATING
C89 m2_2472_13022# VGND 0.831538f $ **FLOATING
C90 m2_3592_15598# VGND 5.94344f $ **FLOATING
C91 m2_2584_17838# VGND 4.71527f $ **FLOATING
C92 m2_2864_23326# VGND 4.89346f $ **FLOATING
C93 m2_3592_27358# VGND 4.41841f $ **FLOATING
C94 m2_2584_29654# VGND 4.17312f $ **FLOATING
C95 m2_2808_33406# VGND 4.18017f $ **FLOATING
C96 m2_3592_35982# VGND 4.2612f $ **FLOATING
C97 m2_3592_39062# VGND 5.95916f $ **FLOATING
C98 m2_3592_42086# VGND 4.35263f $ **FLOATING
C99 vout VGND 98.676704f
C100 clkb VGND 16.841198f
C101 clka VGND 32.197956f
C102 dw_19800_30000# VGND 22.1302f $ **FLOATING
C103 stage1.n0 VGND 0.035278f
C104 stage1.n1 VGND 1.3801f
C105 stage1.t4 VGND 48.4045f
C106 stage1.t0 VGND 0.082135f
C107 stage1.t1 VGND 1.96445f
C108 stage1.t3 VGND 0.079966f
C109 stage1.n2 VGND 0.041838f
C110 stage1.n3 VGND 0.058955f
C111 stage1.n4 VGND 0.058955f
C112 stage1.t2 VGND 1.72035f
C113 stage1.n5 VGND 0.059019f
C114 stage1.n7 VGND 1.03182f
C115 stage1.n8 VGND 0.058955f
C116 stage1.n10 VGND 1.05319f
C117 stage1.n11 VGND 0.045369f
C118 stage1.n12 VGND 0.050911f
C119 stage1.n13 VGND 0.078034f
C120 stage1.n14 VGND 0.169751f
C121 stage1.n15 VGND 0.169751f
C122 stage1.n16 VGND 0.614204f
C123 stage1.n17 VGND 0.078084f
C124 stage1.n18 VGND 0.170037f
C125 stage1.n19 VGND 0.622947f
C126 stage1.n20 VGND 0.614204f
C127 stage1.n21 VGND 0.622947f
C128 stage1.n22 VGND 0.170037f
C129 stage1.n23 VGND 0.06418f
C130 VPWR.t5 VGND 0.003038f
C131 VPWR.n0 VGND 0.007327f
C132 VPWR.t1 VGND 0.003036f
C133 VPWR.n1 VGND 0.003132f
C134 VPWR.n2 VGND 0.003257f
C135 VPWR.n3 VGND 0.003257f
C136 VPWR.n4 VGND 0.003257f
C137 VPWR.t0 VGND 0.052347f
C138 VPWR.n5 VGND 0.003257f
C139 VPWR.n6 VGND 0.003257f
C140 VPWR.n7 VGND 0.00161f
C141 VPWR.n8 VGND 0.003059f
C142 VPWR.n9 VGND 0.003208f
C143 VPWR.n10 VGND 0.003208f
C144 VPWR.n11 VGND 0.040931f
C145 VPWR.n12 VGND 0.003208f
C146 VPWR.n13 VGND 0.003208f
C147 VPWR.n14 VGND 0.003257f
C148 VPWR.n15 VGND 0.001796f
C149 VPWR.n16 VGND 0.003208f
C150 VPWR.n17 VGND 0.040931f
C151 VPWR.n18 VGND 0.003208f
C152 VPWR.n19 VGND 0.001726f
C153 VPWR.n20 VGND 0.001607f
C154 VPWR.n21 VGND 0.004455f
C155 VPWR.n22 VGND 0.012893f
C156 VPWR.t2 VGND 0.385055f
C157 VPWR.t4 VGND 0.015767f
C158 VPWR.n23 VGND 0.140432f
C159 VPWR.n24 VGND 0.008313f
C160 VPWR.n25 VGND 0.011539f
C161 VPWR.n26 VGND 0.011539f
C162 VPWR.t3 VGND 0.33671f
C163 VPWR.n27 VGND 0.011551f
C164 VPWR.n29 VGND 0.201951f
C165 VPWR.n30 VGND 0.011539f
C166 VPWR.n32 VGND 0.206132f
C167 VPWR.n33 VGND 0.008813f
C168 VPWR.n34 VGND 0.006552f
C169 VPWR.n35 VGND 0.009005f
C170 VPWR.n36 VGND 0.01027f
C171 VPWR.n37 VGND 0.015273f
C172 VPWR.n38 VGND 0.033224f
C173 VPWR.n39 VGND 0.033224f
C174 VPWR.n40 VGND 0.120213f
C175 VPWR.n41 VGND 0.015283f
C176 VPWR.n42 VGND 0.03328f
C177 VPWR.n43 VGND 0.121925f
C178 VPWR.n44 VGND 0.120213f
C179 VPWR.n45 VGND 0.121925f
C180 VPWR.n46 VGND 0.03328f
C181 VPWR.n47 VGND 0.012283f
C182 VPWR.n48 VGND 0.009678f
C183 VPWR.n49 VGND 0.129525f
C184 VPWR.n50 VGND 1.41234f
C185 stage3.n0 VGND 0.032636f
C186 stage3.t4 VGND 47.8291f
C187 stage3.t3 VGND 0.077522f
C188 stage3.t0 VGND 1.91766f
C189 stage3.t2 VGND 0.077969f
C190 stage3.n1 VGND 0.044103f
C191 stage3.n2 VGND 0.057545f
C192 stage3.n3 VGND 1.02688f
C193 stage3.n4 VGND 1.00606f
C194 stage3.t1 VGND 0.838692f
C195 stage3.n5 VGND 0.838692f
C196 stage3.n6 VGND 0.057482f
C197 stage3.n7 VGND 0.057482f
C198 stage3.n8 VGND 0.057482f
C199 stage3.n9 VGND 0.041221f
C200 stage3.n10 VGND 0.061605f
C201 stage3.n11 VGND 0.076134f
C202 stage3.n12 VGND 0.16579f
C203 stage3.n13 VGND 0.16579f
C204 stage3.n14 VGND 0.60739f
C205 stage3.n15 VGND 0.076085f
C206 stage3.n16 VGND 0.165511f
C207 stage3.n17 VGND 0.598865f
C208 stage3.n18 VGND 0.60739f
C209 stage3.n19 VGND 0.598865f
C210 stage3.n20 VGND 0.165511f
C211 stage3.n21 VGND 0.050586f
C212 clkb.t2 VGND 58.603302f
C213 clkb.t1 VGND 0.020864f
C214 clkb.t0 VGND 0.032902f
C215 stage2.t3 VGND 1.80979f
C216 stage2.t4 VGND 62.691597f
C217 stage2.t0 VGND 0.096294f
C218 stage2.t1 VGND 2.54782f
C219 stage2.n0 VGND 0.054262f
C220 stage2.n1 VGND 0.076462f
C221 stage2.n2 VGND 0.076462f
C222 stage2.t2 VGND 1.11561f
C223 stage2.n3 VGND 1.11561f
C224 stage2.n4 VGND 0.076546f
C225 stage2.n5 VGND 1.33824f
C226 stage2.n6 VGND 0.076462f
C227 stage2.n7 VGND 1.36594f
C228 stage2.n8 VGND 0.058842f
C229 clka.t2 VGND 0.080865f
C230 clka.t0 VGND 60.1965f
C231 clka.t1 VGND 58.862103f
C232 clka.n0 VGND 2.94109f
.ends

